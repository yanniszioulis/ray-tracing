module pixel_buffer(
    input aclk,
    input aresetn,

    input [7:0] r1, g1, b1,
    input [7:0] r2, g2, b2,
    input [7:0] r3, g3, b3,
    input [7:0] r4, g4, b4,

    input valid1,
    input valid2,
    input valid3,
    input valid4,
    input [2:0] no_of_extra_cores,

    output reg compute_ready_1,
    output reg compute_ready_2,
    output reg compute_ready_3,
    output reg compute_ready_4,

    input in_stream_ready,

    output reg [7:0] out_r,
    output reg [7:0] out_g,
    output reg [7:0] out_b,
    output reg out_valid
);

// State machine states
typedef enum logic [2:0] {
    IDLE,
    WRITE_PIXEL
} state_t;

state_t state, next_state;

// Buffer to store incoming pixels
localparam MAX_CORES = 4;
reg [7:0] pixel_buffer_r[MAX_CORES-1:0];
reg [7:0] pixel_buffer_g[MAX_CORES-1:0];
reg [7:0] pixel_buffer_b[MAX_CORES-1:0];
reg [MAX_CORES-1:0] pixel_buffer_valid;

// Current pixel index to be written next
reg [$clog2(MAX_CORES)-1:0] current_pixel;

// Sequential logic to update state and buffer
always @(posedge aclk or negedge aresetn) begin
    if (!aresetn) begin
        state <= IDLE;
        pixel_buffer_valid <= 'b0;
        current_pixel <= 'b0;
    end else begin
        state <= next_state;

        // Latching valid input pixels into buffer based on the number of enabled cores
        if (valid1 && current_pixel < (no_of_extra_cores + 1)) begin
            pixel_buffer_r[current_pixel] <= r1;
            pixel_buffer_g[current_pixel] <= g1;
            pixel_buffer_b[current_pixel] <= b1;
            pixel_buffer_valid[current_pixel] <= 1'b1;
        end
        if (valid2 && current_pixel < (no_of_extra_cores + 1)) begin
            pixel_buffer_r[current_pixel] <= r2;
            pixel_buffer_g[current_pixel] <= g2;
            pixel_buffer_b[current_pixel] <= b2;
            pixel_buffer_valid[current_pixel] <= 1'b1;
        end
        if (valid3 && current_pixel < (no_of_extra_cores + 1)) begin
            pixel_buffer_r[current_pixel] <= r3;
            pixel_buffer_g[current_pixel] <= g3;
            pixel_buffer_b[current_pixel] <= b3;
            pixel_buffer_valid[current_pixel] <= 1'b1;
        end
        if (valid4 && current_pixel < (no_of_extra_cores + 1)) begin
            pixel_buffer_r[current_pixel] <= r4;
            pixel_buffer_g[current_pixel] <= g4;
            pixel_buffer_b[current_pixel] <= b4;
            pixel_buffer_valid[current_pixel] <= 1'b1;
        end

        // Shifting buffer if pixel is written to packer
        if (state == WRITE_PIXEL && in_stream_ready) begin
            pixel_buffer_valid[current_pixel] <= 1'b0;
            current_pixel <= (current_pixel + 1) % (no_of_extra_cores + 1);
        end
    end
end

// Combinational logic for state transitions and output assignments
always_comb begin
    next_state = state;
    compute_ready_1 = 1'b0;
    compute_ready_2 = 1'b0;
    compute_ready_3 = 1'b0;
    compute_ready_4 = 1'b0;
    out_valid = 1'b0;
    out_r = 8'h00;
    out_g = 8'h00;
    out_b = 8'h00;

    case (state)
        IDLE: begin
            if (pixel_buffer_valid[current_pixel]) begin
                next_state = WRITE_PIXEL;
            end else begin
                case (current_pixel)
                    0: compute_ready_1 = 1'b1;
                    1: compute_ready_2 = 1'b1;
                    2: compute_ready_3 = 1'b1;
                    3: compute_ready_4 = 1'b1;
                endcase
            end
        end

        WRITE_PIXEL: begin
            if (in_stream_ready) begin
                out_r = pixel_buffer_r[current_pixel];
                out_g = pixel_buffer_g[current_pixel];
                out_b = pixel_buffer_b[current_pixel];
                out_valid = 1'b1;
                next_state = IDLE;
            end
        end

        default: begin
            next_state = IDLE;
        end
    endcase
end

endmodule
