module octant_rom #(
    parameter   ADDRESS_WIDTH = 32,
                DATA_WIDTH = 32
)(
    input   logic                       clk,
    input   logic   [ADDRESS_WIDTH-1:0] addr1, addr2,
    output  logic   [DATA_WIDTH-1:0]    dout1, dout2,
    input   logic                       ren1, ren2
);

logic   [DATA_WIDTH-1:0] rom_array [37602:0];

initial begin
    $display("loading mem...");
    $readmemh("effdog.mem", rom_array);
    $display("loaded");
    // rom_array[0] = 32'h00000001;
    // rom_array[1] = 32'h00000009;
    // rom_array[2] = 32'h00000011;
    // rom_array[3] = 32'h00000019;
    // rom_array[4] = 32'h00000021;
    // rom_array[5] = 32'h00000029;
    // rom_array[6] = 32'h00000031;
    // rom_array[7] = 32'h00000039;
    // rom_array[8] = 32'h00000041;
    // rom_array[9] = 32'hFFFFFFF0;
    // rom_array[10] = 32'hFFFFFFF0;
    // rom_array[11] = 32'hFFFFFFF0;
    // rom_array[12] = 32'h00000049;
    // rom_array[13] = 32'hFFFFFFF0;
    // rom_array[14] = 32'hFFFFFFF0;
    // rom_array[15] = 32'hFFFFFFF0;
    // rom_array[16] = 32'h00000051;
    // rom_array[17] = 32'hFFFFFFF0;
    // rom_array[18] = 32'hFFFFFFF0;
    // rom_array[19] = 32'h00000059;
    // rom_array[20] = 32'hFFFFFFF0;
    // rom_array[21] = 32'hFFFFFFF0;
    // rom_array[22] = 32'hFFFFFFF0;
    // rom_array[23] = 32'h00000061;
    // rom_array[24] = 32'hFFFFFFF0;
    // rom_array[25] = 32'hFFFFFFF0;
    // rom_array[26] = 32'h00000069;
    // rom_array[27] = 32'hFFFFFFF0;
    // rom_array[28] = 32'hFFFFFFF0;
    // rom_array[29] = 32'hFFFFFFF0;
    // rom_array[30] = 32'h00000071;
    // rom_array[31] = 32'hFFFFFFF0;
    // rom_array[32] = 32'hFFFFFFF0;
    // rom_array[33] = 32'h00000079;
    // rom_array[34] = 32'hFFFFFFF0;
    // rom_array[35] = 32'hFFFFFFF0;
    // rom_array[36] = 32'hFFFFFFF0;
    // rom_array[37] = 32'h00000081;
    // rom_array[38] = 32'hFFFFFFF0;
    // rom_array[39] = 32'hFFFFFFF0;
    // rom_array[40] = 32'hFFFFFFF0;
    // rom_array[41] = 32'hFFFFFFF0;
    // rom_array[42] = 32'hFFFFFFF0;
    // rom_array[43] = 32'hFFFFFFF0;
    // rom_array[44] = 32'h00000089;
    // rom_array[45] = 32'hFFFFFFF0;
    // rom_array[46] = 32'hFFFFFFF0;
    // rom_array[47] = 32'hFFFFFFF0;
    // rom_array[48] = 32'h00000091;
    // rom_array[49] = 32'hFFFFFFF0;
    // rom_array[50] = 32'hFFFFFFF0;
    // rom_array[51] = 32'h00000099;
    // rom_array[52] = 32'hFFFFFFF0;
    // rom_array[53] = 32'hFFFFFFF0;
    // rom_array[54] = 32'hFFFFFFF0;
    // rom_array[55] = 32'h000000a1;
    // rom_array[56] = 32'hFFFFFFF0;
    // rom_array[57] = 32'hFFFFFFF0;
    // rom_array[58] = 32'h000000a9;
    // rom_array[59] = 32'hFFFFFFF0;
    // rom_array[60] = 32'hFFFFFFF0;
    // rom_array[61] = 32'hFFFFFFF0;
    // rom_array[62] = 32'h000000b1;
    // rom_array[63] = 32'hFFFFFFF0;
    // rom_array[64] = 32'hFFFFFFF0;
    // rom_array[65] = 32'h000000b9;
    // rom_array[66] = 32'hFFFFFFF0;
    // rom_array[67] = 32'hFFFFFFF0;
    // rom_array[68] = 32'hFFFFFFF0;
    // rom_array[69] = 32'h000000c1;
    // rom_array[70] = 32'hFFFFFFF0;
    // rom_array[71] = 32'hFFFFFFF0;
    // rom_array[72] = 32'hFFFFFFF0;
    // rom_array[73] = 32'hFFFFFFF0;
    // rom_array[74] = 32'hFFFFFFF0;
    // rom_array[75] = 32'hFFFFFFF0;
    // rom_array[76] = 32'h000000c9;
    // rom_array[77] = 32'hFFFFFFF0;
    // rom_array[78] = 32'hFFFFFFF0;
    // rom_array[79] = 32'hFFFFFFF0;
    // rom_array[80] = 32'h000000d1;
    // rom_array[81] = 32'hFFFFFFF0;
    // rom_array[82] = 32'hFFFFFFF0;
    // rom_array[83] = 32'hFFFFFFF0;
    // rom_array[84] = 32'h000000d9;
    // rom_array[85] = 32'hFFFFFFF0;
    // rom_array[86] = 32'hFFFFFFF0;
    // rom_array[87] = 32'hFFFFFFF0;
    // rom_array[88] = 32'h000000e1;
    // rom_array[89] = 32'hFFFFFFF0;
    // rom_array[90] = 32'hFFFFFFF0;
    // rom_array[91] = 32'h000000e9;
    // rom_array[92] = 32'hFFFFFFF0;
    // rom_array[93] = 32'hFFFFFFF0;
    // rom_array[94] = 32'hFFFFFFF0;
    // rom_array[95] = 32'h000000f1;
    // rom_array[96] = 32'hFFFFFFF0;
    // rom_array[97] = 32'hFFFFFFF0;
    // rom_array[98] = 32'hFFFFFFF0;
    // rom_array[99] = 32'h000000f9;
    // rom_array[100] = 32'hFFFFFFF0;
    // rom_array[101] = 32'hFFFFFFF0;
    // rom_array[102] = 32'hFFFFFFF0;
    // rom_array[103] = 32'h00000101;
    // rom_array[104] = 32'hFFFFFFF0;
    // rom_array[105] = 32'hFFFFFFF0;
    // rom_array[106] = 32'h00000109;
    // rom_array[107] = 32'hFFFFFFF0;
    // rom_array[108] = 32'hFFFFFFF0;
    // rom_array[109] = 32'hFFFFFFF0;
    // rom_array[110] = 32'h00000111;
    // rom_array[111] = 32'hFFFFFFF0;
    // rom_array[112] = 32'hFFFFFFF0;
    // rom_array[113] = 32'hFFFFFFF0;
    // rom_array[114] = 32'h00000119;
    // rom_array[115] = 32'hFFFFFFF0;
    // rom_array[116] = 32'hFFFFFFF0;
    // rom_array[117] = 32'hFFFFFFF0;
    // rom_array[118] = 32'h00000121;
    // rom_array[119] = 32'hFFFFFFF0;
    // rom_array[120] = 32'hFFFFFFF0;
    // rom_array[121] = 32'h00000129;
    // rom_array[122] = 32'hFFFFFFF0;
    // rom_array[123] = 32'hFFFFFFF0;
    // rom_array[124] = 32'hFFFFFFF0;
    // rom_array[125] = 32'h00000131;
    // rom_array[126] = 32'hFFFFFFF0;
    // rom_array[127] = 32'hFFFFFFF0;
    // rom_array[128] = 32'hFFFFFFF0;
    // rom_array[129] = 32'h00000139;
    // rom_array[130] = 32'hFFFFFFF0;
    // rom_array[131] = 32'hFFFFFFF0;
    // rom_array[132] = 32'hFFFFFFF0;
    // rom_array[133] = 32'h00000141;
    // rom_array[134] = 32'hFFFFFFF0;
    // rom_array[135] = 32'hFFFFFFF0;
    // rom_array[136] = 32'hFFFFFFF0;
    // rom_array[137] = 32'hFFFFFFF0;
    // rom_array[138] = 32'hFFFFFFF0;
    // rom_array[139] = 32'hFFFFFFF0;
    // rom_array[140] = 32'h00000149;
    // rom_array[141] = 32'hFFFFFFF0;
    // rom_array[142] = 32'hFFFFFFF0;
    // rom_array[143] = 32'hFFFFFFF0;
    // rom_array[144] = 32'h00000151;
    // rom_array[145] = 32'hFFFFFFF0;
    // rom_array[146] = 32'hFFFFFFF0;
    // rom_array[147] = 32'hFFFFFFF0;
    // rom_array[148] = 32'h00000159;
    // rom_array[149] = 32'hFFFFFFF0;
    // rom_array[150] = 32'hFFFFFFF0;
    // rom_array[151] = 32'hFFFFFFF0;
    // rom_array[152] = 32'h00000161;
    // rom_array[153] = 32'hFFFFFFF0;
    // rom_array[154] = 32'hFFFFFFF0;
    // rom_array[155] = 32'h00000169;
    // rom_array[156] = 32'hFFFFFFF0;
    // rom_array[157] = 32'hFFFFFFF0;
    // rom_array[158] = 32'hFFFFFFF0;
    // rom_array[159] = 32'h00000171;
    // rom_array[160] = 32'hFFFFFFF0;
    // rom_array[161] = 32'hFFFFFFF0;
    // rom_array[162] = 32'hFFFFFFF0;
    // rom_array[163] = 32'h00000179;
    // rom_array[164] = 32'hFFFFFFF0;
    // rom_array[165] = 32'hFFFFFFF0;
    // rom_array[166] = 32'hFFFFFFF0;
    // rom_array[167] = 32'h00000181;
    // rom_array[168] = 32'hFFFFFFF0;
    // rom_array[169] = 32'hFFFFFFF0;
    // rom_array[170] = 32'h00000189;
    // rom_array[171] = 32'hFFFFFFF0;
    // rom_array[172] = 32'hFFFFFFF0;
    // rom_array[173] = 32'hFFFFFFF0;
    // rom_array[174] = 32'h00000191;
    // rom_array[175] = 32'hFFFFFFF0;
    // rom_array[176] = 32'hFFFFFFF0;
    // rom_array[177] = 32'hFFFFFFF0;
    // rom_array[178] = 32'h00000199;
    // rom_array[179] = 32'hFFFFFFF0;
    // rom_array[180] = 32'hFFFFFFF0;
    // rom_array[181] = 32'hFFFFFFF0;
    // rom_array[182] = 32'hFFFFFFF0;
    // rom_array[183] = 32'hFFFFFFF0;
    // rom_array[184] = 32'hFFFFFFF0;
    // rom_array[185] = 32'h000001a1;
    // rom_array[186] = 32'hFFFFFFF0;
    // rom_array[187] = 32'hFFFFFFF0;
    // rom_array[188] = 32'hFFFFFFF0;
    // rom_array[189] = 32'h000001a9;
    // rom_array[190] = 32'hFFFFFFF0;
    // rom_array[191] = 32'hFFFFFFF0;
    // rom_array[192] = 32'hFFFFFFF0;
    // rom_array[193] = 32'h000001b1;
    // rom_array[194] = 32'hFFFFFFF0;
    // rom_array[195] = 32'hFFFFFFF0;
    // rom_array[196] = 32'hFFFFFFF0;
    // rom_array[197] = 32'hFFFFFFF0;
    // rom_array[198] = 32'hFFFFFFF0;
    // rom_array[199] = 32'hFFFFFFF0;
    // rom_array[200] = 32'hFFFFFFF0;
    // rom_array[201] = 32'hFFFFFFF0;
    // rom_array[202] = 32'hFFFFFFF0;
    // rom_array[203] = 32'hFFFFFFF0;
    // rom_array[204] = 32'hFFFFFFF0;
    // rom_array[205] = 32'hFFFFFFF0;
    // rom_array[206] = 32'hFFFFFFF0;
    // rom_array[207] = 32'hFFFFFFF0;
    // rom_array[208] = 32'h000001b9;
    // rom_array[209] = 32'hFFFFFFF0;
    // rom_array[210] = 32'hFFFFFFF0;
    // rom_array[211] = 32'hFFFFFFF0;
    // rom_array[212] = 32'h000001c1;
    // rom_array[213] = 32'hFFFFFFF0;
    // rom_array[214] = 32'hFFFFFFF0;
    // rom_array[215] = 32'hFFFFFFF0;
    // rom_array[216] = 32'h000001c9;
    // rom_array[217] = 32'hFFFFFFF0;
    // rom_array[218] = 32'hFFFFFFF0;
    // rom_array[219] = 32'hFFFFFFF0;
    // rom_array[220] = 32'h000001d1;
    // rom_array[221] = 32'hFFFFFFF0;
    // rom_array[222] = 32'hFFFFFFF0;
    // rom_array[223] = 32'hFFFFFFF0;
    // rom_array[224] = 32'h000001d9;
    // rom_array[225] = 32'hFFFFFFF0;
    // rom_array[226] = 32'hFFFFFFF0;
    // rom_array[227] = 32'hFFFFFFF0;
    // rom_array[228] = 32'h000001e1;
    // rom_array[229] = 32'hFFFFFFF0;
    // rom_array[230] = 32'hFFFFFFF0;
    // rom_array[231] = 32'hFFFFFFF0;
    // rom_array[232] = 32'h000001e9;
    // rom_array[233] = 32'hFFFFFFF0;
    // rom_array[234] = 32'hFFFFFFF0;
    // rom_array[235] = 32'hFFFFFFF0;
    // rom_array[236] = 32'hFFFFFFF0;
    // rom_array[237] = 32'hFFFFFFF0;
    // rom_array[238] = 32'hFFFFFFF0;
    // rom_array[239] = 32'h000001f1;
    // rom_array[240] = 32'hFFFFFFF0;
    // rom_array[241] = 32'hFFFFFFF0;
    // rom_array[242] = 32'hFFFFFFF0;
    // rom_array[243] = 32'h000001f9;
    // rom_array[244] = 32'hFFFFFFF0;
    // rom_array[245] = 32'hFFFFFFF0;
    // rom_array[246] = 32'hFFFFFFF0;
    // rom_array[247] = 32'h00000201;
    // rom_array[248] = 32'hFFFFFFF0;
    // rom_array[249] = 32'hFFFFFFF0;
    // rom_array[250] = 32'hFFFFFFF0;
    // rom_array[251] = 32'h00000209;
    // rom_array[252] = 32'hFFFFFFF0;
    // rom_array[253] = 32'hFFFFFFF0;
    // rom_array[254] = 32'hFFFFFFF0;
    // rom_array[255] = 32'h00000211;
    // rom_array[256] = 32'hFFFFFFF0;
    // rom_array[257] = 32'hFFFFFFF0;
    // rom_array[258] = 32'hFFFFFFF0;
    // rom_array[259] = 32'h00000219;
    // rom_array[260] = 32'hFFFFFFF0;
    // rom_array[261] = 32'hFFFFFFF0;
    // rom_array[262] = 32'hFFFFFFF0;
    // rom_array[263] = 32'h00000221;
    // rom_array[264] = 32'hFFFFFFF0;
    // rom_array[265] = 32'hFFFFFFF0;
    // rom_array[266] = 32'hFFFFFFF0;
    // rom_array[267] = 32'hFFFFFFF0;
    // rom_array[268] = 32'hFFFFFFF0;
    // rom_array[269] = 32'hFFFFFFF0;
    // rom_array[270] = 32'h00000229;
    // rom_array[271] = 32'hFFFFFFF0;
    // rom_array[272] = 32'hFFFFFFF0;
    // rom_array[273] = 32'hFFFFFFF0;
    // rom_array[274] = 32'h00000231;
    // rom_array[275] = 32'hFFFFFFF0;
    // rom_array[276] = 32'hFFFFFFF0;
    // rom_array[277] = 32'hFFFFFFF0;
    // rom_array[278] = 32'h00000239;
    // rom_array[279] = 32'hFFFFFFF0;
    // rom_array[280] = 32'hFFFFFFF0;
    // rom_array[281] = 32'hFFFFFFF0;
    // rom_array[282] = 32'h00000241;
    // rom_array[283] = 32'hFFFFFFF0;
    // rom_array[284] = 32'hFFFFFFF0;
    // rom_array[285] = 32'hFFFFFFF0;
    // rom_array[286] = 32'h00000249;
    // rom_array[287] = 32'hFFFFFFF0;
    // rom_array[288] = 32'hFFFFFFF0;
    // rom_array[289] = 32'hFFFFFFF0;
    // rom_array[290] = 32'h00000251;
    // rom_array[291] = 32'hFFFFFFF0;
    // rom_array[292] = 32'hFFFFFFF0;
    // rom_array[293] = 32'hFFFFFFF0;
    // rom_array[294] = 32'h00000259;
    // rom_array[295] = 32'hFFFFFFF0;
    // rom_array[296] = 32'hFFFFFFF0;
    // rom_array[297] = 32'hFFFFFFF0;
    // rom_array[298] = 32'hFFFFFFF0;
    // rom_array[299] = 32'hFFFFFFF0;
    // rom_array[300] = 32'hFFFFFFF0;
    // rom_array[301] = 32'h00000261;
    // rom_array[302] = 32'hFFFFFFF0;
    // rom_array[303] = 32'hFFFFFFF0;
    // rom_array[304] = 32'hFFFFFFF0;
    // rom_array[305] = 32'h00000269;
    // rom_array[306] = 32'hFFFFFFF0;
    // rom_array[307] = 32'hFFFFFFF0;
    // rom_array[308] = 32'hFFFFFFF0;
    // rom_array[309] = 32'h00000271;
    // rom_array[310] = 32'hFFFFFFF0;
    // rom_array[311] = 32'hFFFFFFF0;
    // rom_array[312] = 32'hFFFFFFF0;
    // rom_array[313] = 32'h00000279;
    // rom_array[314] = 32'hFFFFFFF0;
    // rom_array[315] = 32'hFFFFFFF0;
    // rom_array[316] = 32'hFFFFFFF0;
    // rom_array[317] = 32'h00000281;
    // rom_array[318] = 32'hFFFFFFF0;
    // rom_array[319] = 32'hFFFFFFF0;
    // rom_array[320] = 32'hFFFFFFF0;
    // rom_array[321] = 32'h00000289;
    // rom_array[322] = 32'hFFFFFFF0;
    // rom_array[323] = 32'hFFFFFFF0;
    // rom_array[324] = 32'hFFFFFFF0;
    // rom_array[325] = 32'h00000291;
    // rom_array[326] = 32'hFFFFFFF0;
    // rom_array[327] = 32'hFFFFFFF0;
    // rom_array[328] = 32'hFFFFFFF0;
    // rom_array[329] = 32'hFFFFFFF0;
    // rom_array[330] = 32'hFFFFFFF0;
    // rom_array[331] = 32'hFFFFFFF0;
    // rom_array[332] = 32'h00000299;
    // rom_array[333] = 32'hFFFFFFF0;
    // rom_array[334] = 32'hFFFFFFF0;
    // rom_array[335] = 32'hFFFFFFF0;
    // rom_array[336] = 32'h000002a1;
    // rom_array[337] = 32'hFFFFFFF0;
    // rom_array[338] = 32'hFFFFFFF0;
    // rom_array[339] = 32'hFFFFFFF0;
    // rom_array[340] = 32'h000002a9;
    // rom_array[341] = 32'hFFFFFFF0;
    // rom_array[342] = 32'hFFFFFFF0;
    // rom_array[343] = 32'hFFFFFFF0;
    // rom_array[344] = 32'h000002b1;
    // rom_array[345] = 32'hFFFFFFF0;
    // rom_array[346] = 32'hFFFFFFF0;
    // rom_array[347] = 32'hFFFFFFF0;
    // rom_array[348] = 32'h000002b9;
    // rom_array[349] = 32'hFFFFFFF0;
    // rom_array[350] = 32'hFFFFFFF0;
    // rom_array[351] = 32'hFFFFFFF0;
    // rom_array[352] = 32'h000002c1;
    // rom_array[353] = 32'hFFFFFFF0;
    // rom_array[354] = 32'hFFFFFFF0;
    // rom_array[355] = 32'hFFFFFFF0;
    // rom_array[356] = 32'h000002c9;
    // rom_array[357] = 32'hFFFFFFF0;
    // rom_array[358] = 32'hFFFFFFF0;
    // rom_array[359] = 32'hFFFFFFF0;
    // rom_array[360] = 32'hFFFFFFF0;
    // rom_array[361] = 32'hFFFFFFF0;
    // rom_array[362] = 32'hFFFFFFF0;
    // rom_array[363] = 32'h000002d1;
    // rom_array[364] = 32'hFFFFFFF0;
    // rom_array[365] = 32'hFFFFFFF0;
    // rom_array[366] = 32'hFFFFFFF0;
    // rom_array[367] = 32'h000002d9;
    // rom_array[368] = 32'hFFFFFFF0;
    // rom_array[369] = 32'hFFFFFFF0;
    // rom_array[370] = 32'hFFFFFFF0;
    // rom_array[371] = 32'h000002e1;
    // rom_array[372] = 32'hFFFFFFF0;
    // rom_array[373] = 32'hFFFFFFF0;
    // rom_array[374] = 32'hFFFFFFF0;
    // rom_array[375] = 32'h000002e9;
    // rom_array[376] = 32'hFFFFFFF0;
    // rom_array[377] = 32'hFFFFFFF0;
    // rom_array[378] = 32'hFFFFFFF0;
    // rom_array[379] = 32'h000002f1;
    // rom_array[380] = 32'hFFFFFFF0;
    // rom_array[381] = 32'hFFFFFFF0;
    // rom_array[382] = 32'hFFFFFFF0;
    // rom_array[383] = 32'h000002f9;
    // rom_array[384] = 32'hFFFFFFF0;
    // rom_array[385] = 32'hFFFFFFF0;
    // rom_array[386] = 32'hFFFFFFF0;
    // rom_array[387] = 32'h00000301;
    // rom_array[388] = 32'hFFFFFFF0;
    // rom_array[389] = 32'hFFFFFFF0;
    // rom_array[390] = 32'hFFFFFFF0;
    // rom_array[391] = 32'hFFFFFFF0;
    // rom_array[392] = 32'hFFFFFFF0;
    // rom_array[393] = 32'hFFFFFFF0;
    // rom_array[394] = 32'h00000309;
    // rom_array[395] = 32'hFFFFFFF0;
    // rom_array[396] = 32'hFFFFFFF0;
    // rom_array[397] = 32'hFFFFFFF0;
    // rom_array[398] = 32'h00000311;
    // rom_array[399] = 32'hFFFFFFF0;
    // rom_array[400] = 32'hFFFFFFF0;
    // rom_array[401] = 32'hFFFFFFF0;
    // rom_array[402] = 32'h00000319;
    // rom_array[403] = 32'hFFFFFFF0;
    // rom_array[404] = 32'hFFFFFFF0;
    // rom_array[405] = 32'hFFFFFFF0;
    // rom_array[406] = 32'h00000321;
    // rom_array[407] = 32'hFFFFFFF0;
    // rom_array[408] = 32'hFFFFFFF0;
    // rom_array[409] = 32'hFFFFFFF0;
    // rom_array[410] = 32'h00000329;
    // rom_array[411] = 32'hFFFFFFF0;
    // rom_array[412] = 32'hFFFFFFF0;
    // rom_array[413] = 32'hFFFFFFF0;
    // rom_array[414] = 32'h00000331;
    // rom_array[415] = 32'hFFFFFFF0;
    // rom_array[416] = 32'hFFFFFFF0;
    // rom_array[417] = 32'h00000339;
    // rom_array[418] = 32'hFFFFFFF0;
    // rom_array[419] = 32'hFFFFFFF0;
    // rom_array[420] = 32'hFFFFFFF0;
    // rom_array[421] = 32'h00000341;
    // rom_array[422] = 32'hFFFFFFF0;
    // rom_array[423] = 32'hFFFFFFF0;
    // rom_array[424] = 32'hFFFFFFF0;
    // rom_array[425] = 32'h00000349;
    // rom_array[426] = 32'hFFFFFFF0;
    // rom_array[427] = 32'hFFFFFFF0;
    // rom_array[428] = 32'hFFFFFFF0;
    // rom_array[429] = 32'h00000351;
    // rom_array[430] = 32'hFFFFFFF0;
    // rom_array[431] = 32'hFFFFFFF0;
    // rom_array[432] = 32'hFFFFFFF0;
    // rom_array[433] = 32'h00000359;
    // rom_array[434] = 32'hFFFFFFF0;
    // rom_array[435] = 32'hFFFFFFF0;
    // rom_array[436] = 32'hFFFFFFF0;
    // rom_array[437] = 32'h00000361;
    // rom_array[438] = 32'hFFFFFFF0;
    // rom_array[439] = 32'hFFFFFFF0;
    // rom_array[440] = 32'hFFFFFFF0;
    // rom_array[441] = 32'hFFFFFFF0;
    // rom_array[442] = 32'hFFFFFFF0;
    // rom_array[443] = 32'hFFFFFFF0;
    // rom_array[444] = 32'hFFFFFFF0;
    // rom_array[445] = 32'hFFFFFFF0;
    // rom_array[446] = 32'h00000369;
    // rom_array[447] = 32'hFFFFFFF0;
    // rom_array[448] = 32'h00000371;
    // rom_array[449] = 32'hFFFFFFF0;
    // rom_array[450] = 32'h00000379;
    // rom_array[451] = 32'hFFFFFFF0;
    // rom_array[452] = 32'h00000381;
    // rom_array[453] = 32'hFFFFFFF0;
    // rom_array[454] = 32'h00000389;
    // rom_array[455] = 32'hFFFFFFF0;
    // rom_array[456] = 32'h00000391;
    // rom_array[457] = 32'hFFFFFFF0;
    // rom_array[458] = 32'h00000399;
    // rom_array[459] = 32'hFFFFFFF0;
    // rom_array[460] = 32'h000003a1;
    // rom_array[461] = 32'hFFFFFFF0;
    // rom_array[462] = 32'h000003a9;
    // rom_array[463] = 32'hFFFFFFF0;
    // rom_array[464] = 32'h000003b1;
    // rom_array[465] = 32'hFFFFFFF0;
    // rom_array[466] = 32'hFFFFFFF0;
    // rom_array[467] = 32'hFFFFFFF0;
    // rom_array[468] = 32'h000003b9;
    // rom_array[469] = 32'hFFFFFFF0;
    // rom_array[470] = 32'h000003c1;
    // rom_array[471] = 32'hFFFFFFF0;
    // rom_array[472] = 32'h000003c9;
    // rom_array[473] = 32'hFFFFFFF0;
    // rom_array[474] = 32'hFFFFFFF0;
    // rom_array[475] = 32'hFFFFFFF0;
    // rom_array[476] = 32'hFFFFFFF0;
    // rom_array[477] = 32'hFFFFFFF0;
    // rom_array[478] = 32'h000003d1;
    // rom_array[479] = 32'hFFFFFFF0;
    // rom_array[480] = 32'h000003d9;
    // rom_array[481] = 32'hFFFFFFF0;
    // rom_array[482] = 32'hFFFFFFF0;
    // rom_array[483] = 32'hFFFFFFF0;
    // rom_array[484] = 32'h000003e1;
    // rom_array[485] = 32'hFFFFFFF0;
    // rom_array[486] = 32'hFFFFFFF0;
    // rom_array[487] = 32'hFFFFFFF0;
    // rom_array[488] = 32'hFFFFFFF0;
    // rom_array[489] = 32'hFFFFFFF0;
    // rom_array[490] = 32'h000003e9;
    // rom_array[491] = 32'hFFFFFFF0;
    // rom_array[492] = 32'h000003f1;
    // rom_array[493] = 32'hFFFFFFF0;
    // rom_array[494] = 32'h000003f9;
    // rom_array[495] = 32'hFFFFFFF0;
    // rom_array[496] = 32'h00000401;
    // rom_array[497] = 32'hFFFFFFF0;
    // rom_array[498] = 32'hFFFFFFF0;
    // rom_array[499] = 32'hFFFFFFF0;
    // rom_array[500] = 32'hFFFFFFF0;
    // rom_array[501] = 32'h00000409;
    // rom_array[502] = 32'hFFFFFFF0;
    // rom_array[503] = 32'h00000411;
    // rom_array[504] = 32'hFFFFFFF0;
    // rom_array[505] = 32'h00000419;
    // rom_array[506] = 32'hFFFFFFF0;
    // rom_array[507] = 32'h00000421;
    // rom_array[508] = 32'hFFFFFFF0;
    // rom_array[509] = 32'h00000429;
    // rom_array[510] = 32'hFFFFFFF0;
    // rom_array[511] = 32'h00000431;
    // rom_array[512] = 32'hFFFFFFF0;
    // rom_array[513] = 32'h00000439;
    // rom_array[514] = 32'hFFFFFFF0;
    // rom_array[515] = 32'h00000441;
    // rom_array[516] = 32'hFFFFFFF0;
    // rom_array[517] = 32'h00000449;
    // rom_array[518] = 32'hFFFFFFF0;
    // rom_array[519] = 32'h00000451;
    // rom_array[520] = 32'hFFFFFFF0;
    // rom_array[521] = 32'hFFFFFFF0;
    // rom_array[522] = 32'hFFFFFFF0;
    // rom_array[523] = 32'h00000459;
    // rom_array[524] = 32'hFFFFFFF0;
    // rom_array[525] = 32'h00000461;
    // rom_array[526] = 32'hFFFFFFF0;
    // rom_array[527] = 32'h00000469;
    // rom_array[528] = 32'hFFFFFFF0;
    // rom_array[529] = 32'hFFFFFFF0;
    // rom_array[530] = 32'hFFFFFFF0;
    // rom_array[531] = 32'hFFFFFFF0;
    // rom_array[532] = 32'hFFFFFFF0;
    // rom_array[533] = 32'h00000471;
    // rom_array[534] = 32'hFFFFFFF0;
    // rom_array[535] = 32'h00000479;
    // rom_array[536] = 32'hFFFFFFF0;
    // rom_array[537] = 32'hFFFFFFF0;
    // rom_array[538] = 32'hFFFFFFF0;
    // rom_array[539] = 32'h00000481;
    // rom_array[540] = 32'hFFFFFFF0;
    // rom_array[541] = 32'hFFFFFFF0;
    // rom_array[542] = 32'hFFFFFFF0;
    // rom_array[543] = 32'hFFFFFFF0;
    // rom_array[544] = 32'hFFFFFFF0;
    // rom_array[545] = 32'h00000489;
    // rom_array[546] = 32'hFFFFFFF0;
    // rom_array[547] = 32'h00000491;
    // rom_array[548] = 32'hFFFFFFF0;
    // rom_array[549] = 32'h00000499;
    // rom_array[550] = 32'hFFFFFFF0;
    // rom_array[551] = 32'h000004a1;
    // rom_array[552] = 32'hFFFFFFF0;
    // rom_array[553] = 32'hFFFFFFF0;
    // rom_array[554] = 32'hFFFFFFF0;
    // rom_array[555] = 32'hFFFFFFF0;
    // rom_array[556] = 32'hFFFFFFF0;
    // rom_array[557] = 32'hFFFFFFF0;
    // rom_array[558] = 32'h000004a9;
    // rom_array[559] = 32'hFFFFFFF0;
    // rom_array[560] = 32'h000004b1;
    // rom_array[561] = 32'hFFFFFFF0;
    // rom_array[562] = 32'h000004b9;
    // rom_array[563] = 32'hFFFFFFF0;
    // rom_array[564] = 32'h000004c1;
    // rom_array[565] = 32'hFFFFFFF0;
    // rom_array[566] = 32'h000004c9;
    // rom_array[567] = 32'hFFFFFFF0;
    // rom_array[568] = 32'h000004d1;
    // rom_array[569] = 32'hFFFFFFF0;
    // rom_array[570] = 32'h000004d9;
    // rom_array[571] = 32'hFFFFFFF0;
    // rom_array[572] = 32'h000004e1;
    // rom_array[573] = 32'hFFFFFFF0;
    // rom_array[574] = 32'h000004e9;
    // rom_array[575] = 32'hFFFFFFF0;
    // rom_array[576] = 32'h000004f1;
    // rom_array[577] = 32'hFFFFFFF0;
    // rom_array[578] = 32'h000004f9;
    // rom_array[579] = 32'hFFFFFFF0;
    // rom_array[580] = 32'h00000501;
    // rom_array[581] = 32'hFFFFFFF0;
    // rom_array[582] = 32'h00000509;
    // rom_array[583] = 32'hFFFFFFF0;
    // rom_array[584] = 32'h00000511;
    // rom_array[585] = 32'hFFFFFFF0;
    // rom_array[586] = 32'hFFFFFFF0;
    // rom_array[587] = 32'hFFFFFFF0;
    // rom_array[588] = 32'hFFFFFFF0;
    // rom_array[589] = 32'hFFFFFFF0;
    // rom_array[590] = 32'h00000519;
    // rom_array[591] = 32'hFFFFFFF0;
    // rom_array[592] = 32'h00000521;
    // rom_array[593] = 32'hFFFFFFF0;
    // rom_array[594] = 32'h00000529;
    // rom_array[595] = 32'hFFFFFFF0;
    // rom_array[596] = 32'h00000531;
    // rom_array[597] = 32'hFFFFFFF0;
    // rom_array[598] = 32'hFFFFFFF0;
    // rom_array[599] = 32'hFFFFFFF0;
    // rom_array[600] = 32'hFFFFFFF0;
    // rom_array[601] = 32'hFFFFFFF0;
    // rom_array[602] = 32'h00000539;
    // rom_array[603] = 32'hFFFFFFF0;
    // rom_array[604] = 32'h00000541;
    // rom_array[605] = 32'hFFFFFFF0;
    // rom_array[606] = 32'h00000549;
    // rom_array[607] = 32'hFFFFFFF0;
    // rom_array[608] = 32'h00000551;
    // rom_array[609] = 32'hFFFFFFF0;
    // rom_array[610] = 32'hFFFFFFF0;
    // rom_array[611] = 32'hFFFFFFF0;
    // rom_array[612] = 32'hFFFFFFF0;
    // rom_array[613] = 32'h00000559;
    // rom_array[614] = 32'hFFFFFFF0;
    // rom_array[615] = 32'h00000561;
    // rom_array[616] = 32'hFFFFFFF0;
    // rom_array[617] = 32'h00000569;
    // rom_array[618] = 32'hFFFFFFF0;
    // rom_array[619] = 32'h00000571;
    // rom_array[620] = 32'hFFFFFFF0;
    // rom_array[621] = 32'h00000579;
    // rom_array[622] = 32'hFFFFFFF0;
    // rom_array[623] = 32'h00000581;
    // rom_array[624] = 32'hFFFFFFF0;
    // rom_array[625] = 32'h00000589;
    // rom_array[626] = 32'hFFFFFFF0;
    // rom_array[627] = 32'h00000591;
    // rom_array[628] = 32'hFFFFFFF0;
    // rom_array[629] = 32'h00000599;
    // rom_array[630] = 32'hFFFFFFF0;
    // rom_array[631] = 32'h000005a1;
    // rom_array[632] = 32'hFFFFFFF0;
    // rom_array[633] = 32'h000005a9;
    // rom_array[634] = 32'hFFFFFFF0;
    // rom_array[635] = 32'h000005b1;
    // rom_array[636] = 32'hFFFFFFF0;
    // rom_array[637] = 32'h000005b9;
    // rom_array[638] = 32'hFFFFFFF0;
    // rom_array[639] = 32'h000005c1;
    // rom_array[640] = 32'hFFFFFFF0;
    // rom_array[641] = 32'hFFFFFFF0;
    // rom_array[642] = 32'hFFFFFFF0;
    // rom_array[643] = 32'hFFFFFFF0;
    // rom_array[644] = 32'hFFFFFFF0;
    // rom_array[645] = 32'h000005c9;
    // rom_array[646] = 32'hFFFFFFF0;
    // rom_array[647] = 32'h000005d1;
    // rom_array[648] = 32'hFFFFFFF0;
    // rom_array[649] = 32'h000005d9;
    // rom_array[650] = 32'hFFFFFFF0;
    // rom_array[651] = 32'h000005e1;
    // rom_array[652] = 32'hFFFFFFF0;
    // rom_array[653] = 32'hFFFFFFF0;
    // rom_array[654] = 32'hFFFFFFF0;
    // rom_array[655] = 32'hFFFFFFF0;
    // rom_array[656] = 32'hFFFFFFF0;
    // rom_array[657] = 32'h000005e9;
    // rom_array[658] = 32'hFFFFFFF0;
    // rom_array[659] = 32'h000005f1;
    // rom_array[660] = 32'hFFFFFFF0;
    // rom_array[661] = 32'h000005f9;
    // rom_array[662] = 32'hFFFFFFF0;
    // rom_array[663] = 32'h00000601;
    // rom_array[664] = 32'hFFFFFFF0;
    // rom_array[665] = 32'hFFFFFFF0;
    // rom_array[666] = 32'h00000609;
    // rom_array[667] = 32'hFFFFFFF0;
    // rom_array[668] = 32'h00000611;
    // rom_array[669] = 32'hFFFFFFF0;
    // rom_array[670] = 32'h00000619;
    // rom_array[671] = 32'hFFFFFFF0;
    // rom_array[672] = 32'h00000621;
    // rom_array[673] = 32'hFFFFFFF0;
    // rom_array[674] = 32'h00000629;
    // rom_array[675] = 32'hFFFFFFF0;
    // rom_array[676] = 32'h00000631;
    // rom_array[677] = 32'hFFFFFFF0;
    // rom_array[678] = 32'h00000639;
    // rom_array[679] = 32'hFFFFFFF0;
    // rom_array[680] = 32'h00000641;
    // rom_array[681] = 32'hFFFFFFF0;
    // rom_array[682] = 32'h00000649;
    // rom_array[683] = 32'hFFFFFFF0;
    // rom_array[684] = 32'h00000651;
    // rom_array[685] = 32'hFFFFFFF0;
    // rom_array[686] = 32'h00000659;
    // rom_array[687] = 32'hFFFFFFF0;
    // rom_array[688] = 32'h00000661;
    // rom_array[689] = 32'hFFFFFFF0;
    // rom_array[690] = 32'hFFFFFFF0;
    // rom_array[691] = 32'hFFFFFFF0;
    // rom_array[692] = 32'hFFFFFFF0;
    // rom_array[693] = 32'hFFFFFFF0;
    // rom_array[694] = 32'h00000669;
    // rom_array[695] = 32'hFFFFFFF0;
    // rom_array[696] = 32'h00000671;
    // rom_array[697] = 32'hFFFFFFF0;
    // rom_array[698] = 32'h00000679;
    // rom_array[699] = 32'hFFFFFFF0;
    // rom_array[700] = 32'h00000681;
    // rom_array[701] = 32'hFFFFFFF0;
    // rom_array[702] = 32'h00000689;
    // rom_array[703] = 32'hFFFFFFF0;
    // rom_array[704] = 32'h00000691;
    // rom_array[705] = 32'hFFFFFFF0;
    // rom_array[706] = 32'h00000699;
    // rom_array[707] = 32'hFFFFFFF0;
    // rom_array[708] = 32'h000006a1;
    // rom_array[709] = 32'hFFFFFFF0;
    // rom_array[710] = 32'h000006a9;
    // rom_array[711] = 32'hFFFFFFF0;
    // rom_array[712] = 32'h000006b1;
    // rom_array[713] = 32'hFFFFFFF0;
    // rom_array[714] = 32'h000006b9;
    // rom_array[715] = 32'hFFFFFFF0;
    // rom_array[716] = 32'h000006c1;
    // rom_array[717] = 32'hFFFFFFF0;
    // rom_array[718] = 32'hFFFFFFF0;
    // rom_array[719] = 32'hFFFFFFF0;
    // rom_array[720] = 32'hFFFFFFF0;
    // rom_array[721] = 32'h000006c9;
    // rom_array[722] = 32'hFFFFFFF0;
    // rom_array[723] = 32'h000006d1;
    // rom_array[724] = 32'hFFFFFFF0;
    // rom_array[725] = 32'h000006d9;
    // rom_array[726] = 32'hFFFFFFF0;
    // rom_array[727] = 32'h000006e1;
    // rom_array[728] = 32'hFFFFFFF0;
    // rom_array[729] = 32'h000006e9;
    // rom_array[730] = 32'hFFFFFFF0;
    // rom_array[731] = 32'h000006f1;
    // rom_array[732] = 32'hFFFFFFF0;
    // rom_array[733] = 32'h000006f9;
    // rom_array[734] = 32'hFFFFFFF0;
    // rom_array[735] = 32'h00000701;
    // rom_array[736] = 32'hFFFFFFF0;
    // rom_array[737] = 32'h00000709;
    // rom_array[738] = 32'hFFFFFFF0;
    // rom_array[739] = 32'h00000711;
    // rom_array[740] = 32'hFFFFFFF0;
    // rom_array[741] = 32'h00000719;
    // rom_array[742] = 32'hFFFFFFF0;
    // rom_array[743] = 32'h00000721;
    // rom_array[744] = 32'hFFFFFFF0;
    // rom_array[745] = 32'hFFFFFFF0;
    // rom_array[746] = 32'hFFFFFFF0;
    // rom_array[747] = 32'hFFFFFFF0;
    // rom_array[748] = 32'hFFFFFFF0;
    // rom_array[749] = 32'h00000729;
    // rom_array[750] = 32'hFFFFFFF0;
    // rom_array[751] = 32'h00000731;
    // rom_array[752] = 32'hFFFFFFF0;
    // rom_array[753] = 32'h00000739;
    // rom_array[754] = 32'hFFFFFFF0;
    // rom_array[755] = 32'h00000741;
    // rom_array[756] = 32'hFFFFFFF0;
    // rom_array[757] = 32'h00000749;
    // rom_array[758] = 32'hFFFFFFF0;
    // rom_array[759] = 32'h00000751;
    // rom_array[760] = 32'hFFFFFFF0;
    // rom_array[761] = 32'h00000759;
    // rom_array[762] = 32'hFFFFFFF0;
    // rom_array[763] = 32'h00000761;
    // rom_array[764] = 32'hFFFFFFF0;
    // rom_array[765] = 32'h00000769;
    // rom_array[766] = 32'hFFFFFFF0;
    // rom_array[767] = 32'h00000771;
    // rom_array[768] = 32'hFFFFFFF0;
    // rom_array[769] = 32'h00000779;
    // rom_array[770] = 32'hFFFFFFF0;
    // rom_array[771] = 32'h00000781;
    // rom_array[772] = 32'hFFFFFFF0;
    // rom_array[773] = 32'hFFFFFFF0;
    // rom_array[774] = 32'hFFFFFFF0;
    // rom_array[775] = 32'hFFFFFFF0;
    // rom_array[776] = 32'hFFFFFFF0;
    // rom_array[777] = 32'hFFFFFFF0;
    // rom_array[778] = 32'h00000789;
    // rom_array[779] = 32'hFFFFFFF0;
    // rom_array[780] = 32'h00000791;
    // rom_array[781] = 32'hFFFFFFF0;
    // rom_array[782] = 32'h00000799;
    // rom_array[783] = 32'hFFFFFFF0;
    // rom_array[784] = 32'h000007a1;
    // rom_array[785] = 32'hFFFFFFF0;
    // rom_array[786] = 32'h000007a9;
    // rom_array[787] = 32'hFFFFFFF0;
    // rom_array[788] = 32'h000007b1;
    // rom_array[789] = 32'hFFFFFFF0;
    // rom_array[790] = 32'h000007b9;
    // rom_array[791] = 32'hFFFFFFF0;
    // rom_array[792] = 32'hFFFFFFF0;
    // rom_array[793] = 32'hFFFFFFF0;
    // rom_array[794] = 32'h000007c1;
    // rom_array[795] = 32'hFFFFFFF0;
    // rom_array[796] = 32'h000007c9;
    // rom_array[797] = 32'hFFFFFFF0;
    // rom_array[798] = 32'h000007d1;
    // rom_array[799] = 32'hFFFFFFF0;
    // rom_array[800] = 32'h000007d9;
    // rom_array[801] = 32'hFFFFFFF0;
    // rom_array[802] = 32'hFFFFFFF0;
    // rom_array[803] = 32'hFFFFFFF0;
    // rom_array[804] = 32'hFFFFFFF0;
    // rom_array[805] = 32'hFFFFFFF0;
    // rom_array[806] = 32'h000007e1;
    // rom_array[807] = 32'hFFFFFFF0;
    // rom_array[808] = 32'h000007e9;
    // rom_array[809] = 32'hFFFFFFF0;
    // rom_array[810] = 32'h000007f1;
    // rom_array[811] = 32'hFFFFFFF0;
    // rom_array[812] = 32'h000007f9;
    // rom_array[813] = 32'hFFFFFFF0;
    // rom_array[814] = 32'h00000801;
    // rom_array[815] = 32'hFFFFFFF0;
    // rom_array[816] = 32'h00000809;
    // rom_array[817] = 32'hFFFFFFF0;
    // rom_array[818] = 32'h00000811;
    // rom_array[819] = 32'hFFFFFFF0;
    // rom_array[820] = 32'h00000819;
    // rom_array[821] = 32'hFFFFFFF0;
    // rom_array[822] = 32'h00000821;
    // rom_array[823] = 32'hFFFFFFF0;
    // rom_array[824] = 32'h00000829;
    // rom_array[825] = 32'h00000831;
    // rom_array[826] = 32'hFFFFFFF0;
    // rom_array[827] = 32'h00000839;
    // rom_array[828] = 32'hFFFFFFF0;
    // rom_array[829] = 32'h00000841;
    // rom_array[830] = 32'hFFFFFFF0;
    // rom_array[831] = 32'h00000849;
    // rom_array[832] = 32'hFFFFFFF0;
    // rom_array[833] = 32'h00000851;
    // rom_array[834] = 32'hFFFFFFF0;
    // rom_array[835] = 32'h00000859;
    // rom_array[836] = 32'hFFFFFFF0;
    // rom_array[837] = 32'h00000861;
    // rom_array[838] = 32'hFFFFFFF0;
    // rom_array[839] = 32'hFFFFFFF0;
    // rom_array[840] = 32'hFFFFFFF0;
    // rom_array[841] = 32'h00000869;
    // rom_array[842] = 32'hFFFFFFF0;
    // rom_array[843] = 32'h00000871;
    // rom_array[844] = 32'hFFFFFFF0;
    // rom_array[845] = 32'h00000879;
    // rom_array[846] = 32'hFFFFFFF0;
    // rom_array[847] = 32'h00000881;
    // rom_array[848] = 32'hFFFFFFF0;
    // rom_array[849] = 32'hFFFFFFF0;
    // rom_array[850] = 32'hFFFFFFF0;
    // rom_array[851] = 32'hFFFFFFF0;
    // rom_array[852] = 32'hFFFFFFF0;
    // rom_array[853] = 32'h00000889;
    // rom_array[854] = 32'hFFFFFFF0;
    // rom_array[855] = 32'h00000891;
    // rom_array[856] = 32'hFFFFFFF0;
    // rom_array[857] = 32'h00000899;
    // rom_array[858] = 32'hFFFFFFF0;
    // rom_array[859] = 32'h000008a1;
    // rom_array[860] = 32'hFFFFFFF0;
    // rom_array[861] = 32'h000008a9;
    // rom_array[862] = 32'hFFFFFFF0;
    // rom_array[863] = 32'h000008b1;
    // rom_array[864] = 32'hFFFFFFF0;
    // rom_array[865] = 32'h000008b9;
    // rom_array[866] = 32'hFFFFFFF0;
    // rom_array[867] = 32'h000008c1;
    // rom_array[868] = 32'hFFFFFFF0;
    // rom_array[869] = 32'h000008c9;
    // rom_array[870] = 32'hFFFFFFF0;
    // rom_array[871] = 32'h000008d1;
    // rom_array[872] = 32'hFFFFFFF0;
    // rom_array[873] = 32'hFFFFFFF0;
    // rom_array[874] = 32'hFFFFFFF0;
    // rom_array[875] = 32'hFFFFFFF0;
    // rom_array[876] = 32'hFFFFFFF0;
    // rom_array[877] = 32'hFFFFFFF0;
    // rom_array[878] = 32'hFFFFFFF0;
    // rom_array[879] = 32'hFFFFFFF0;
    // rom_array[880] = 32'h000008d9;
    // rom_array[881] = 32'hFFFFFFF0;
    // rom_array[882] = 32'hFFFFFFF0;
    // rom_array[883] = 32'hFFFFFFF0;
    // rom_array[884] = 32'hFFFFFFF0;
    // rom_array[885] = 32'hFFFFFFF0;
    // rom_array[886] = 32'h000008e1;
    // rom_array[887] = 32'hFFFFFFF0;
    // rom_array[888] = 32'hFFFFFFF0;
    // rom_array[889] = 32'hFFFFFFF0;
    // rom_array[890] = 32'hFFFFFFF0;
    // rom_array[891] = 32'hFFFFFFF0;
    // rom_array[892] = 32'h000008e9;
    // rom_array[893] = 32'hFFFFFFF0;
    // rom_array[894] = 32'hFFFFFFF0;
    // rom_array[895] = 32'hFFFFFFF0;
    // rom_array[896] = 32'h000008f1;
    // rom_array[897] = 32'hFFFFFFF0;
    // rom_array[898] = 32'h000008f9;
    // rom_array[899] = 32'hFFFFFFF0;
    // rom_array[900] = 32'h00000901;
    // rom_array[901] = 32'hFFFFFFF0;
    // rom_array[902] = 32'h00000909;
    // rom_array[903] = 32'hFFFFFFF0;
    // rom_array[904] = 32'h00000911;
    // rom_array[905] = 32'hFFFFFFF0;
    // rom_array[906] = 32'hFFFFFFF0;
    // rom_array[907] = 32'hFFFFFFF0;
    // rom_array[908] = 32'h00000919;
    // rom_array[909] = 32'hFFFFFFF0;
    // rom_array[910] = 32'hFFFFFFF0;
    // rom_array[911] = 32'hFFFFFFF0;
    // rom_array[912] = 32'hFFFFFFF0;
    // rom_array[913] = 32'hFFFFFFF0;
    // rom_array[914] = 32'h00000921;
    // rom_array[915] = 32'hFFFFFFF0;
    // rom_array[916] = 32'hFFFFFFF0;
    // rom_array[917] = 32'hFFFFFFF0;
    // rom_array[918] = 32'hFFFFFFF0;
    // rom_array[919] = 32'hFFFFFFF0;
    // rom_array[920] = 32'hFFFFFFF0;
    // rom_array[921] = 32'hFFFFFFF0;
    // rom_array[922] = 32'hFFFFFFF0;
    // rom_array[923] = 32'hFFFFFFF0;
    // rom_array[924] = 32'hFFFFFFF0;
    // rom_array[925] = 32'hFFFFFFF0;
    // rom_array[926] = 32'hFFFFFFF0;
    // rom_array[927] = 32'hFFFFFFF0;
    // rom_array[928] = 32'h00000929;
    // rom_array[929] = 32'hFFFFFFF0;
    // rom_array[930] = 32'hFFFFFFF0;
    // rom_array[931] = 32'hFFFFFFF0;
    // rom_array[932] = 32'hFFFFFFF0;
    // rom_array[933] = 32'hFFFFFFF0;
    // rom_array[934] = 32'h00000931;
    // rom_array[935] = 32'hFFFFFFF0;
    // rom_array[936] = 32'h00000939;
    // rom_array[937] = 32'hFFFFFFF0;
    // rom_array[938] = 32'hFFFFFFF0;
    // rom_array[939] = 32'hFFFFFFF0;
    // rom_array[940] = 32'h00000941;
    // rom_array[941] = 32'hFFFFFFF0;
    // rom_array[942] = 32'hFFFFFFF0;
    // rom_array[943] = 32'hFFFFFFF0;
    // rom_array[944] = 32'hFFFFFFF0;
    // rom_array[945] = 32'hFFFFFFF0;
    // rom_array[946] = 32'h00000949;
    // rom_array[947] = 32'hFFFFFFF0;
    // rom_array[948] = 32'h00000951;
    // rom_array[949] = 32'hFFFFFFF0;
    // rom_array[950] = 32'h00000959;
    // rom_array[951] = 32'hFFFFFFF0;
    // rom_array[952] = 32'h00000961;
    // rom_array[953] = 32'hFFFFFFF0;
    // rom_array[954] = 32'h00000969;
    // rom_array[955] = 32'hFFFFFFF0;
    // rom_array[956] = 32'h00000971;
    // rom_array[957] = 32'hFFFFFFF0;
    // rom_array[958] = 32'h00000979;
    // rom_array[959] = 32'hFFFFFFF0;
    // rom_array[960] = 32'h00000981;
    // rom_array[961] = 32'hFFFFFFF0;
    // rom_array[962] = 32'hFFFFFFF0;
    // rom_array[963] = 32'hFFFFFFF0;
    // rom_array[964] = 32'h00000989;
    // rom_array[965] = 32'hFFFFFFF0;
    // rom_array[966] = 32'hFFFFFFF0;
    // rom_array[967] = 32'hFFFFFFF0;
    // rom_array[968] = 32'h00000991;
    // rom_array[969] = 32'hFFFFFFF0;
    // rom_array[970] = 32'h00000999;
    // rom_array[971] = 32'hFFFFFFF0;
    // rom_array[972] = 32'h000009a1;
    // rom_array[973] = 32'hFFFFFFF0;
    // rom_array[974] = 32'h000009a9;
    // rom_array[975] = 32'hFFFFFFF0;
    // rom_array[976] = 32'h000009b1;
    // rom_array[977] = 32'hFFFFFFF0;
    // rom_array[978] = 32'hFFFFFFF0;
    // rom_array[979] = 32'hFFFFFFF0;
    // rom_array[980] = 32'h000009b9;
    // rom_array[981] = 32'hFFFFFFF0;
    // rom_array[982] = 32'hFFFFFFF0;
    // rom_array[983] = 32'hFFFFFFF0;
    // rom_array[984] = 32'h000009c1;
    // rom_array[985] = 32'hFFFFFFF0;
    // rom_array[986] = 32'h000009c9;
    // rom_array[987] = 32'hFFFFFFF0;
    // rom_array[988] = 32'h000009d1;
    // rom_array[989] = 32'hFFFFFFF0;
    // rom_array[990] = 32'h000009d9;
    // rom_array[991] = 32'hFFFFFFF0;
    // rom_array[992] = 32'h000009e1;
    // rom_array[993] = 32'hFFFFFFF0;
    // rom_array[994] = 32'hFFFFFFF0;
    // rom_array[995] = 32'hFFFFFFF0;
    // rom_array[996] = 32'h000009e9;
    // rom_array[997] = 32'hFFFFFFF0;
    // rom_array[998] = 32'hFFFFFFF0;
    // rom_array[999] = 32'hFFFFFFF0;
    // rom_array[1000] = 32'h000009f1;
    // rom_array[1001] = 32'hFFFFFFF0;
    // rom_array[1002] = 32'hFFFFFFF0;
    // rom_array[1003] = 32'hFFFFFFF0;
    // rom_array[1004] = 32'h000009f9;
    // rom_array[1005] = 32'hFFFFFFF0;
    // rom_array[1006] = 32'hFFFFFFF0;
    // rom_array[1007] = 32'hFFFFFFF0;
    // rom_array[1008] = 32'h00000a01;
    // rom_array[1009] = 32'hFFFFFFF0;
    // rom_array[1010] = 32'h00000a09;
    // rom_array[1011] = 32'hFFFFFFF0;
    // rom_array[1012] = 32'h00000a11;
    // rom_array[1013] = 32'hFFFFFFF0;
    // rom_array[1014] = 32'h00000a19;
    // rom_array[1015] = 32'hFFFFFFF0;
    // rom_array[1016] = 32'h00000a21;
    // rom_array[1017] = 32'hFFFFFFF0;
    // rom_array[1018] = 32'hFFFFFFF0;
    // rom_array[1019] = 32'hFFFFFFF0;
    // rom_array[1020] = 32'h00000a29;
    // rom_array[1021] = 32'hFFFFFFF0;
    // rom_array[1022] = 32'hFFFFFFF0;
    // rom_array[1023] = 32'hFFFFFFF0;
    // rom_array[1024] = 32'h00000a31;
    // rom_array[1025] = 32'hFFFFFFF0;
    // rom_array[1026] = 32'h00000a39;
    // rom_array[1027] = 32'hFFFFFFF0;
    // rom_array[1028] = 32'h00000a41;
    // rom_array[1029] = 32'hFFFFFFF0;
    // rom_array[1030] = 32'h00000a49;
    // rom_array[1031] = 32'hFFFFFFF0;
    // rom_array[1032] = 32'h00000a51;
    // rom_array[1033] = 32'hFFFFFFF0;
    // rom_array[1034] = 32'hFFFFFFF0;
    // rom_array[1035] = 32'hFFFFFFF0;
    // rom_array[1036] = 32'hFFFFFFF0;
    // rom_array[1037] = 32'hFFFFFFF0;
    // rom_array[1038] = 32'hFFFFFFF0;
    // rom_array[1039] = 32'h00000a59;
    // rom_array[1040] = 32'hFFFFFFF0;
    // rom_array[1041] = 32'hFFFFFFF0;
    // rom_array[1042] = 32'hFFFFFFF0;
    // rom_array[1043] = 32'hFFFFFFF0;
    // rom_array[1044] = 32'hFFFFFFF0;
    // rom_array[1045] = 32'h00000a61;
    // rom_array[1046] = 32'hFFFFFFF0;
    // rom_array[1047] = 32'hFFFFFFF0;
    // rom_array[1048] = 32'hFFFFFFF0;
    // rom_array[1049] = 32'hFFFFFFF0;
    // rom_array[1050] = 32'hFFFFFFF0;
    // rom_array[1051] = 32'h00000a69;
    // rom_array[1052] = 32'hFFFFFFF0;
    // rom_array[1053] = 32'hFFFFFFF0;
    // rom_array[1054] = 32'hFFFFFFF0;
    // rom_array[1055] = 32'h00000a71;
    // rom_array[1056] = 32'hFFFFFFF0;
    // rom_array[1057] = 32'h00000a79;
    // rom_array[1058] = 32'hFFFFFFF0;
    // rom_array[1059] = 32'h00000a81;
    // rom_array[1060] = 32'hFFFFFFF0;
    // rom_array[1061] = 32'h00000a89;
    // rom_array[1062] = 32'hFFFFFFF0;
    // rom_array[1063] = 32'h00000a91;
    // rom_array[1064] = 32'hFFFFFFF0;
    // rom_array[1065] = 32'hFFFFFFF0;
    // rom_array[1066] = 32'hFFFFFFF0;
    // rom_array[1067] = 32'h00000a99;
    // rom_array[1068] = 32'hFFFFFFF0;
    // rom_array[1069] = 32'hFFFFFFF0;
    // rom_array[1070] = 32'hFFFFFFF0;
    // rom_array[1071] = 32'hFFFFFFF0;
    // rom_array[1072] = 32'hFFFFFFF0;
    // rom_array[1073] = 32'h00000aa1;
    // rom_array[1074] = 32'hFFFFFFF0;
    // rom_array[1075] = 32'hFFFFFFF0;
    // rom_array[1076] = 32'hFFFFFFF0;
    // rom_array[1077] = 32'hFFFFFFF0;
    // rom_array[1078] = 32'hFFFFFFF0;
    // rom_array[1079] = 32'hFFFFFFF0;
    // rom_array[1080] = 32'hFFFFFFF0;
    // rom_array[1081] = 32'hFFFFFFF0;
    // rom_array[1082] = 32'hFFFFFFF0;
    // rom_array[1083] = 32'hFFFFFFF0;
    // rom_array[1084] = 32'hFFFFFFF0;
    // rom_array[1085] = 32'hFFFFFFF0;
    // rom_array[1086] = 32'hFFFFFFF0;
    // rom_array[1087] = 32'h00000aa9;
    // rom_array[1088] = 32'hFFFFFFF0;
    // rom_array[1089] = 32'hFFFFFFF0;
    // rom_array[1090] = 32'hFFFFFFF0;
    // rom_array[1091] = 32'hFFFFFFF0;
    // rom_array[1092] = 32'hFFFFFFF0;
    // rom_array[1093] = 32'h00000ab1;
    // rom_array[1094] = 32'hFFFFFFF0;
    // rom_array[1095] = 32'h00000ab9;
    // rom_array[1096] = 32'hFFFFFFF0;
    // rom_array[1097] = 32'hFFFFFFF0;
    // rom_array[1098] = 32'hFFFFFFF0;
    // rom_array[1099] = 32'h00000ac1;
    // rom_array[1100] = 32'hFFFFFFF0;
    // rom_array[1101] = 32'hFFFFFFF0;
    // rom_array[1102] = 32'hFFFFFFF0;
    // rom_array[1103] = 32'hFFFFFFF0;
    // rom_array[1104] = 32'hFFFFFFF0;
    // rom_array[1105] = 32'h00000ac9;
    // rom_array[1106] = 32'hFFFFFFF0;
    // rom_array[1107] = 32'h00000ad1;
    // rom_array[1108] = 32'hFFFFFFF0;
    // rom_array[1109] = 32'h00000ad9;
    // rom_array[1110] = 32'hFFFFFFF0;
    // rom_array[1111] = 32'h00000ae1;
    // rom_array[1112] = 32'hFFFFFFF0;
    // rom_array[1113] = 32'h00000ae9;
    // rom_array[1114] = 32'hFFFFFFF0;
    // rom_array[1115] = 32'h00000af1;
    // rom_array[1116] = 32'hFFFFFFF0;
    // rom_array[1117] = 32'h00000af9;
    // rom_array[1118] = 32'hFFFFFFF0;
    // rom_array[1119] = 32'h00000b01;
    // rom_array[1120] = 32'hFFFFFFF0;
    // rom_array[1121] = 32'hFFFFFFF0;
    // rom_array[1122] = 32'hFFFFFFF0;
    // rom_array[1123] = 32'h00000b09;
    // rom_array[1124] = 32'hFFFFFFF0;
    // rom_array[1125] = 32'hFFFFFFF0;
    // rom_array[1126] = 32'hFFFFFFF0;
    // rom_array[1127] = 32'h00000b11;
    // rom_array[1128] = 32'hFFFFFFF0;
    // rom_array[1129] = 32'h00000b19;
    // rom_array[1130] = 32'hFFFFFFF0;
    // rom_array[1131] = 32'h00000b21;
    // rom_array[1132] = 32'hFFFFFFF0;
    // rom_array[1133] = 32'h00000b29;
    // rom_array[1134] = 32'hFFFFFFF0;
    // rom_array[1135] = 32'h00000b31;
    // rom_array[1136] = 32'hFFFFFFF0;
    // rom_array[1137] = 32'hFFFFFFF0;
    // rom_array[1138] = 32'hFFFFFFF0;
    // rom_array[1139] = 32'h00000b39;
    // rom_array[1140] = 32'hFFFFFFF0;
    // rom_array[1141] = 32'hFFFFFFF0;
    // rom_array[1142] = 32'hFFFFFFF0;
    // rom_array[1143] = 32'h00000b41;
    // rom_array[1144] = 32'hFFFFFFF0;
    // rom_array[1145] = 32'h00000b49;
    // rom_array[1146] = 32'hFFFFFFF0;
    // rom_array[1147] = 32'h00000b51;
    // rom_array[1148] = 32'hFFFFFFF0;
    // rom_array[1149] = 32'h00000b59;
    // rom_array[1150] = 32'hFFFFFFF0;
    // rom_array[1151] = 32'h00000b61;
    // rom_array[1152] = 32'hFFFFFFF0;
    // rom_array[1153] = 32'hFFFFFFF0;
    // rom_array[1154] = 32'hFFFFFFF0;
    // rom_array[1155] = 32'h00000b69;
    // rom_array[1156] = 32'hFFFFFFF0;
    // rom_array[1157] = 32'hFFFFFFF0;
    // rom_array[1158] = 32'hFFFFFFF0;
    // rom_array[1159] = 32'h00000b71;
    // rom_array[1160] = 32'hFFFFFFF0;
    // rom_array[1161] = 32'hFFFFFFF0;
    // rom_array[1162] = 32'hFFFFFFF0;
    // rom_array[1163] = 32'h00000b79;
    // rom_array[1164] = 32'hFFFFFFF0;
    // rom_array[1165] = 32'hFFFFFFF0;
    // rom_array[1166] = 32'hFFFFFFF0;
    // rom_array[1167] = 32'h00000b81;
    // rom_array[1168] = 32'hFFFFFFF0;
    // rom_array[1169] = 32'h00000b89;
    // rom_array[1170] = 32'hFFFFFFF0;
    // rom_array[1171] = 32'h00000b91;
    // rom_array[1172] = 32'hFFFFFFF0;
    // rom_array[1173] = 32'h00000b99;
    // rom_array[1174] = 32'hFFFFFFF0;
    // rom_array[1175] = 32'h00000ba1;
    // rom_array[1176] = 32'hFFFFFFF0;
    // rom_array[1177] = 32'hFFFFFFF0;
    // rom_array[1178] = 32'hFFFFFFF0;
    // rom_array[1179] = 32'h00000ba9;
    // rom_array[1180] = 32'hFFFFFFF0;
    // rom_array[1181] = 32'hFFFFFFF0;
    // rom_array[1182] = 32'hFFFFFFF0;
    // rom_array[1183] = 32'h00000bb1;
    // rom_array[1184] = 32'hFFFFFFF0;
    // rom_array[1185] = 32'h00000bb9;
    // rom_array[1186] = 32'hFFFFFFF0;
    // rom_array[1187] = 32'h00000bc1;
    // rom_array[1188] = 32'hFFFFFFF0;
    // rom_array[1189] = 32'h00000bc9;
    // rom_array[1190] = 32'hFFFFFFF0;
    // rom_array[1191] = 32'h00000bd1;
    // rom_array[1192] = 32'hFFFFFFF0;
    // rom_array[1193] = 32'hFFFFFFF0;
    // rom_array[1194] = 32'hFFFFFFF0;
    // rom_array[1195] = 32'hFFFFFFF0;
    // rom_array[1196] = 32'hFFFFFFF0;
    // rom_array[1197] = 32'hFFFFFFF0;
    // rom_array[1198] = 32'hFFFFFFF0;
    // rom_array[1199] = 32'hFFFFFFF0;
    // rom_array[1200] = 32'h00000bd9;
    // rom_array[1201] = 32'hFFFFFFF0;
    // rom_array[1202] = 32'hFFFFFFF0;
    // rom_array[1203] = 32'hFFFFFFF0;
    // rom_array[1204] = 32'hFFFFFFF0;
    // rom_array[1205] = 32'hFFFFFFF0;
    // rom_array[1206] = 32'h00000be1;
    // rom_array[1207] = 32'hFFFFFFF0;
    // rom_array[1208] = 32'hFFFFFFF0;
    // rom_array[1209] = 32'hFFFFFFF0;
    // rom_array[1210] = 32'h00000be9;
    // rom_array[1211] = 32'hFFFFFFF0;
    // rom_array[1212] = 32'h00000bf1;
    // rom_array[1213] = 32'hFFFFFFF0;
    // rom_array[1214] = 32'h00000bf9;
    // rom_array[1215] = 32'hFFFFFFF0;
    // rom_array[1216] = 32'h00000c01;
    // rom_array[1217] = 32'hFFFFFFF0;
    // rom_array[1218] = 32'h00000c09;
    // rom_array[1219] = 32'hFFFFFFF0;
    // rom_array[1220] = 32'hFFFFFFF0;
    // rom_array[1221] = 32'hFFFFFFF0;
    // rom_array[1222] = 32'h00000c11;
    // rom_array[1223] = 32'hFFFFFFF0;
    // rom_array[1224] = 32'hFFFFFFF0;
    // rom_array[1225] = 32'hFFFFFFF0;
    // rom_array[1226] = 32'hFFFFFFF0;
    // rom_array[1227] = 32'hFFFFFFF0;
    // rom_array[1228] = 32'h00000c19;
    // rom_array[1229] = 32'hFFFFFFF0;
    // rom_array[1230] = 32'hFFFFFFF0;
    // rom_array[1231] = 32'hFFFFFFF0;
    // rom_array[1232] = 32'hFFFFFFF0;
    // rom_array[1233] = 32'hFFFFFFF0;
    // rom_array[1234] = 32'h00000c21;
    // rom_array[1235] = 32'hFFFFFFF0;
    // rom_array[1236] = 32'hFFFFFFF0;
    // rom_array[1237] = 32'hFFFFFFF0;
    // rom_array[1238] = 32'hFFFFFFF0;
    // rom_array[1239] = 32'hFFFFFFF0;
    // rom_array[1240] = 32'hFFFFFFF0;
    // rom_array[1241] = 32'hFFFFFFF0;
    // rom_array[1242] = 32'hFFFFFFF0;
    // rom_array[1243] = 32'hFFFFFFF0;
    // rom_array[1244] = 32'hFFFFFFF0;
    // rom_array[1245] = 32'hFFFFFFF0;
    // rom_array[1246] = 32'h00000c29;
    // rom_array[1247] = 32'hFFFFFFF0;
    // rom_array[1248] = 32'h00000c31;
    // rom_array[1249] = 32'hFFFFFFF0;
    // rom_array[1250] = 32'hFFFFFFF0;
    // rom_array[1251] = 32'hFFFFFFF0;
    // rom_array[1252] = 32'hFFFFFFF0;
    // rom_array[1253] = 32'hFFFFFFF0;
    // rom_array[1254] = 32'h00000c39;
    // rom_array[1255] = 32'hFFFFFFF0;
    // rom_array[1256] = 32'hFFFFFFF0;
    // rom_array[1257] = 32'hFFFFFFF0;
    // rom_array[1258] = 32'h00000c41;
    // rom_array[1259] = 32'hFFFFFFF0;
    // rom_array[1260] = 32'h00000c49;
    // rom_array[1261] = 32'hFFFFFFF0;
    // rom_array[1262] = 32'h00000c51;
    // rom_array[1263] = 32'hFFFFFFF0;
    // rom_array[1264] = 32'h00000c59;
    // rom_array[1265] = 32'hFFFFFFF0;
    // rom_array[1266] = 32'h00000c61;
    // rom_array[1267] = 32'hFFFFFFF0;
    // rom_array[1268] = 32'hFFFFFFF0;
    // rom_array[1269] = 32'hFFFFFFF0;
    // rom_array[1270] = 32'h00000c69;
    // rom_array[1271] = 32'hFFFFFFF0;
    // rom_array[1272] = 32'hFFFFFFF0;
    // rom_array[1273] = 32'hFFFFFFF0;
    // rom_array[1274] = 32'h00000c71;
    // rom_array[1275] = 32'hFFFFFFF0;
    // rom_array[1276] = 32'h00000c79;
    // rom_array[1277] = 32'hFFFFFFF0;
    // rom_array[1278] = 32'h00000c81;
    // rom_array[1279] = 32'hFFFFFFF0;
    // rom_array[1280] = 32'h00000c89;
    // rom_array[1281] = 32'hFFFFFFF0;
    // rom_array[1282] = 32'h00000c91;
    // rom_array[1283] = 32'hFFFFFFF0;
    // rom_array[1284] = 32'hFFFFFFF0;
    // rom_array[1285] = 32'hFFFFFFF0;
    // rom_array[1286] = 32'h00000c99;
    // rom_array[1287] = 32'hFFFFFFF0;
    // rom_array[1288] = 32'hFFFFFFF0;
    // rom_array[1289] = 32'hFFFFFFF0;
    // rom_array[1290] = 32'h00000ca1;
    // rom_array[1291] = 32'hFFFFFFF0;
    // rom_array[1292] = 32'h00000ca9;
    // rom_array[1293] = 32'hFFFFFFF0;
    // rom_array[1294] = 32'h00000cb1;
    // rom_array[1295] = 32'hFFFFFFF0;
    // rom_array[1296] = 32'h00000cb9;
    // rom_array[1297] = 32'hFFFFFFF0;
    // rom_array[1298] = 32'h00000cc1;
    // rom_array[1299] = 32'hFFFFFFF0;
    // rom_array[1300] = 32'hFFFFFFF0;
    // rom_array[1301] = 32'hFFFFFFF0;
    // rom_array[1302] = 32'h00000cc9;
    // rom_array[1303] = 32'hFFFFFFF0;
    // rom_array[1304] = 32'hFFFFFFF0;
    // rom_array[1305] = 32'hFFFFFFF0;
    // rom_array[1306] = 32'h00000cd1;
    // rom_array[1307] = 32'hFFFFFFF0;
    // rom_array[1308] = 32'h00000cd9;
    // rom_array[1309] = 32'hFFFFFFF0;
    // rom_array[1310] = 32'h00000ce1;
    // rom_array[1311] = 32'hFFFFFFF0;
    // rom_array[1312] = 32'h00000ce9;
    // rom_array[1313] = 32'hFFFFFFF0;
    // rom_array[1314] = 32'h00000cf1;
    // rom_array[1315] = 32'hFFFFFFF0;
    // rom_array[1316] = 32'hFFFFFFF0;
    // rom_array[1317] = 32'hFFFFFFF0;
    // rom_array[1318] = 32'h00000cf9;
    // rom_array[1319] = 32'hFFFFFFF0;
    // rom_array[1320] = 32'hFFFFFFF0;
    // rom_array[1321] = 32'hFFFFFFF0;
    // rom_array[1322] = 32'h00000d01;
    // rom_array[1323] = 32'hFFFFFFF0;
    // rom_array[1324] = 32'h00000d09;
    // rom_array[1325] = 32'hFFFFFFF0;
    // rom_array[1326] = 32'h00000d11;
    // rom_array[1327] = 32'hFFFFFFF0;
    // rom_array[1328] = 32'h00000d19;
    // rom_array[1329] = 32'hFFFFFFF0;
    // rom_array[1330] = 32'h00000d21;
    // rom_array[1331] = 32'hFFFFFFF0;
    // rom_array[1332] = 32'hFFFFFFF0;
    // rom_array[1333] = 32'hFFFFFFF0;
    // rom_array[1334] = 32'h00000d29;
    // rom_array[1335] = 32'hFFFFFFF0;
    // rom_array[1336] = 32'hFFFFFFF0;
    // rom_array[1337] = 32'hFFFFFFF0;
    // rom_array[1338] = 32'h00000d31;
    // rom_array[1339] = 32'hFFFFFFF0;
    // rom_array[1340] = 32'h00000d39;
    // rom_array[1341] = 32'hFFFFFFF0;
    // rom_array[1342] = 32'h00000d41;
    // rom_array[1343] = 32'hFFFFFFF0;
    // rom_array[1344] = 32'h00000d49;
    // rom_array[1345] = 32'hFFFFFFF0;
    // rom_array[1346] = 32'h00000d51;
    // rom_array[1347] = 32'hFFFFFFF0;
    // rom_array[1348] = 32'hFFFFFFF0;
    // rom_array[1349] = 32'hFFFFFFF0;
    // rom_array[1350] = 32'h00000d59;
    // rom_array[1351] = 32'hFFFFFFF0;
    // rom_array[1352] = 32'hFFFFFFF0;
    // rom_array[1353] = 32'hFFFFFFF0;
    // rom_array[1354] = 32'h00000d61;
    // rom_array[1355] = 32'hFFFFFFF0;
    // rom_array[1356] = 32'h00000d69;
    // rom_array[1357] = 32'hFFFFFFF0;
    // rom_array[1358] = 32'h00000d71;
    // rom_array[1359] = 32'hFFFFFFF0;
    // rom_array[1360] = 32'h00000d79;
    // rom_array[1361] = 32'hFFFFFFF0;
    // rom_array[1362] = 32'h00000d81;
    // rom_array[1363] = 32'hFFFFFFF0;
    // rom_array[1364] = 32'hFFFFFFF0;
    // rom_array[1365] = 32'hFFFFFFF0;
    // rom_array[1366] = 32'h00000d89;
    // rom_array[1367] = 32'hFFFFFFF0;
    // rom_array[1368] = 32'hFFFFFFF0;
    // rom_array[1369] = 32'hFFFFFFF0;
    // rom_array[1370] = 32'hFFFFFFF0;
    // rom_array[1371] = 32'hFFFFFFF0;
    // rom_array[1372] = 32'hFFFFFFF0;
    // rom_array[1373] = 32'hFFFFFFF0;
    // rom_array[1374] = 32'hFFFFFFF0;
    // rom_array[1375] = 32'h00000d91;
    // rom_array[1376] = 32'hFFFFFFF0;
    // rom_array[1377] = 32'hFFFFFFF0;
    // rom_array[1378] = 32'hFFFFFFF0;
    // rom_array[1379] = 32'hFFFFFFF0;
    // rom_array[1380] = 32'hFFFFFFF0;
    // rom_array[1381] = 32'h00000d99;
    // rom_array[1382] = 32'hFFFFFFF0;
    // rom_array[1383] = 32'hFFFFFFF0;
    // rom_array[1384] = 32'hFFFFFFF0;
    // rom_array[1385] = 32'h00000da1;
    // rom_array[1386] = 32'hFFFFFFF0;
    // rom_array[1387] = 32'h00000da9;
    // rom_array[1388] = 32'hFFFFFFF0;
    // rom_array[1389] = 32'h00000db1;
    // rom_array[1390] = 32'hFFFFFFF0;
    // rom_array[1391] = 32'h00000db9;
    // rom_array[1392] = 32'hFFFFFFF0;
    // rom_array[1393] = 32'h00000dc1;
    // rom_array[1394] = 32'hFFFFFFF0;
    // rom_array[1395] = 32'hFFFFFFF0;
    // rom_array[1396] = 32'hFFFFFFF0;
    // rom_array[1397] = 32'h00000dc9;
    // rom_array[1398] = 32'hFFFFFFF0;
    // rom_array[1399] = 32'hFFFFFFF0;
    // rom_array[1400] = 32'hFFFFFFF0;
    // rom_array[1401] = 32'hFFFFFFF0;
    // rom_array[1402] = 32'hFFFFFFF0;
    // rom_array[1403] = 32'h00000dd1;
    // rom_array[1404] = 32'hFFFFFFF0;
    // rom_array[1405] = 32'hFFFFFFF0;
    // rom_array[1406] = 32'hFFFFFFF0;
    // rom_array[1407] = 32'hFFFFFFF0;
    // rom_array[1408] = 32'hFFFFFFF0;
    // rom_array[1409] = 32'h00000dd9;
    // rom_array[1410] = 32'hFFFFFFF0;
    // rom_array[1411] = 32'hFFFFFFF0;
    // rom_array[1412] = 32'hFFFFFFF0;
    // rom_array[1413] = 32'hFFFFFFF0;
    // rom_array[1414] = 32'hFFFFFFF0;
    // rom_array[1415] = 32'hFFFFFFF0;
    // rom_array[1416] = 32'hFFFFFFF0;
    // rom_array[1417] = 32'hFFFFFFF0;
    // rom_array[1418] = 32'hFFFFFFF0;
    // rom_array[1419] = 32'hFFFFFFF0;
    // rom_array[1420] = 32'hFFFFFFF0;
    // rom_array[1421] = 32'h00000de1;
    // rom_array[1422] = 32'hFFFFFFF0;
    // rom_array[1423] = 32'h00000de9;
    // rom_array[1424] = 32'hFFFFFFF0;
    // rom_array[1425] = 32'hFFFFFFF0;
    // rom_array[1426] = 32'hFFFFFFF0;
    // rom_array[1427] = 32'hFFFFFFF0;
    // rom_array[1428] = 32'hFFFFFFF0;
    // rom_array[1429] = 32'h00000df1;
    // rom_array[1430] = 32'hFFFFFFF0;
    // rom_array[1431] = 32'hFFFFFFF0;
    // rom_array[1432] = 32'hFFFFFFF0;
    // rom_array[1433] = 32'h00000df9;
    // rom_array[1434] = 32'hFFFFFFF0;
    // rom_array[1435] = 32'h00000e01;
    // rom_array[1436] = 32'hFFFFFFF0;
    // rom_array[1437] = 32'h00000e09;
    // rom_array[1438] = 32'hFFFFFFF0;
    // rom_array[1439] = 32'h00000e11;
    // rom_array[1440] = 32'hFFFFFFF0;
    // rom_array[1441] = 32'h00000e19;
    // rom_array[1442] = 32'hFFFFFFF0;
    // rom_array[1443] = 32'hFFFFFFF0;
    // rom_array[1444] = 32'hFFFFFFF0;
    // rom_array[1445] = 32'h00000e21;
    // rom_array[1446] = 32'hFFFFFFF0;
    // rom_array[1447] = 32'hFFFFFFF0;
    // rom_array[1448] = 32'hFFFFFFF0;
    // rom_array[1449] = 32'h00000e29;
    // rom_array[1450] = 32'hFFFFFFF0;
    // rom_array[1451] = 32'h00000e31;
    // rom_array[1452] = 32'hFFFFFFF0;
    // rom_array[1453] = 32'h00000e39;
    // rom_array[1454] = 32'hFFFFFFF0;
    // rom_array[1455] = 32'h00000e41;
    // rom_array[1456] = 32'hFFFFFFF0;
    // rom_array[1457] = 32'h00000e49;
    // rom_array[1458] = 32'hFFFFFFF0;
    // rom_array[1459] = 32'hFFFFFFF0;
    // rom_array[1460] = 32'hFFFFFFF0;
    // rom_array[1461] = 32'h00000e51;
    // rom_array[1462] = 32'hFFFFFFF0;
    // rom_array[1463] = 32'hFFFFFFF0;
    // rom_array[1464] = 32'hFFFFFFF0;
    // rom_array[1465] = 32'h00000e59;
    // rom_array[1466] = 32'hFFFFFFF0;
    // rom_array[1467] = 32'h00000e61;
    // rom_array[1468] = 32'hFFFFFFF0;
    // rom_array[1469] = 32'h00000e69;
    // rom_array[1470] = 32'hFFFFFFF0;
    // rom_array[1471] = 32'h00000e71;
    // rom_array[1472] = 32'hFFFFFFF0;
    // rom_array[1473] = 32'h00000e79;
    // rom_array[1474] = 32'hFFFFFFF0;
    // rom_array[1475] = 32'hFFFFFFF0;
    // rom_array[1476] = 32'hFFFFFFF0;
    // rom_array[1477] = 32'h00000e81;
    // rom_array[1478] = 32'hFFFFFFF0;
    // rom_array[1479] = 32'hFFFFFFF0;
    // rom_array[1480] = 32'hFFFFFFF0;
    // rom_array[1481] = 32'h00000e89;
    // rom_array[1482] = 32'hFFFFFFF0;
    // rom_array[1483] = 32'h00000e91;
    // rom_array[1484] = 32'hFFFFFFF0;
    // rom_array[1485] = 32'h00000e99;
    // rom_array[1486] = 32'hFFFFFFF0;
    // rom_array[1487] = 32'h00000ea1;
    // rom_array[1488] = 32'hFFFFFFF0;
    // rom_array[1489] = 32'h00000ea9;
    // rom_array[1490] = 32'hFFFFFFF0;
    // rom_array[1491] = 32'hFFFFFFF0;
    // rom_array[1492] = 32'hFFFFFFF0;
    // rom_array[1493] = 32'h00000eb1;
    // rom_array[1494] = 32'hFFFFFFF0;
    // rom_array[1495] = 32'hFFFFFFF0;
    // rom_array[1496] = 32'hFFFFFFF0;
    // rom_array[1497] = 32'h00000eb9;
    // rom_array[1498] = 32'hFFFFFFF0;
    // rom_array[1499] = 32'h00000ec1;
    // rom_array[1500] = 32'hFFFFFFF0;
    // rom_array[1501] = 32'h00000ec9;
    // rom_array[1502] = 32'hFFFFFFF0;
    // rom_array[1503] = 32'h00000ed1;
    // rom_array[1504] = 32'hFFFFFFF0;
    // rom_array[1505] = 32'h00000ed9;
    // rom_array[1506] = 32'hFFFFFFF0;
    // rom_array[1507] = 32'hFFFFFFF0;
    // rom_array[1508] = 32'hFFFFFFF0;
    // rom_array[1509] = 32'h00000ee1;
    // rom_array[1510] = 32'hFFFFFFF0;
    // rom_array[1511] = 32'hFFFFFFF0;
    // rom_array[1512] = 32'hFFFFFFF0;
    // rom_array[1513] = 32'h00000ee9;
    // rom_array[1514] = 32'hFFFFFFF0;
    // rom_array[1515] = 32'h00000ef1;
    // rom_array[1516] = 32'hFFFFFFF0;
    // rom_array[1517] = 32'h00000ef9;
    // rom_array[1518] = 32'hFFFFFFF0;
    // rom_array[1519] = 32'h00000f01;
    // rom_array[1520] = 32'hFFFFFFF0;
    // rom_array[1521] = 32'h00000f09;
    // rom_array[1522] = 32'hFFFFFFF0;
    // rom_array[1523] = 32'hFFFFFFF0;
    // rom_array[1524] = 32'hFFFFFFF0;
    // rom_array[1525] = 32'h00000f11;
    // rom_array[1526] = 32'hFFFFFFF0;
    // rom_array[1527] = 32'hFFFFFFF0;
    // rom_array[1528] = 32'hFFFFFFF0;
    // rom_array[1529] = 32'h00000f19;
    // rom_array[1530] = 32'hFFFFFFF0;
    // rom_array[1531] = 32'h00000f21;
    // rom_array[1532] = 32'hFFFFFFF0;
    // rom_array[1533] = 32'h00000f29;
    // rom_array[1534] = 32'hFFFFFFF0;
    // rom_array[1535] = 32'h00000f31;
    // rom_array[1536] = 32'hFFFFFFF0;
    // rom_array[1537] = 32'h00000f39;
    // rom_array[1538] = 32'hFFFFFFF0;
    // rom_array[1539] = 32'hFFFFFFF0;
    // rom_array[1540] = 32'hFFFFFFF0;
    // rom_array[1541] = 32'h00000f41;
    // rom_array[1542] = 32'hFFFFFFF0;
    // rom_array[1543] = 32'hFFFFFFF0;
    // rom_array[1544] = 32'hFFFFFFF0;
    // rom_array[1545] = 32'hFFFFFFF0;
    // rom_array[1546] = 32'hFFFFFFF0;
    // rom_array[1547] = 32'hFFFFFFF0;
    // rom_array[1548] = 32'h00000f49;
    // rom_array[1549] = 32'hFFFFFFF0;
    // rom_array[1550] = 32'hFFFFFFF0;
    // rom_array[1551] = 32'hFFFFFFF0;
    // rom_array[1552] = 32'hFFFFFFF0;
    // rom_array[1553] = 32'hFFFFFFF0;
    // rom_array[1554] = 32'h00000f51;
    // rom_array[1555] = 32'hFFFFFFF0;
    // rom_array[1556] = 32'h00000f59;
    // rom_array[1557] = 32'hFFFFFFF0;
    // rom_array[1558] = 32'hFFFFFFF0;
    // rom_array[1559] = 32'hFFFFFFF0;
    // rom_array[1560] = 32'hFFFFFFF0;
    // rom_array[1561] = 32'hFFFFFFF0;
    // rom_array[1562] = 32'hFFFFFFF0;
    // rom_array[1563] = 32'hFFFFFFF0;
    // rom_array[1564] = 32'h00000f61;
    // rom_array[1565] = 32'hFFFFFFF0;
    // rom_array[1566] = 32'hFFFFFFF0;
    // rom_array[1567] = 32'hFFFFFFF0;
    // rom_array[1568] = 32'h00000f69;
    // rom_array[1569] = 32'hFFFFFFF0;
    // rom_array[1570] = 32'h00000f71;
    // rom_array[1571] = 32'hFFFFFFF0;
    // rom_array[1572] = 32'h00000f79;
    // rom_array[1573] = 32'hFFFFFFF0;
    // rom_array[1574] = 32'h00000f81;
    // rom_array[1575] = 32'hFFFFFFF0;
    // rom_array[1576] = 32'h00000f89;
    // rom_array[1577] = 32'hFFFFFFF0;
    // rom_array[1578] = 32'hFFFFFFF0;
    // rom_array[1579] = 32'hFFFFFFF0;
    // rom_array[1580] = 32'h00000f91;
    // rom_array[1581] = 32'hFFFFFFF0;
    // rom_array[1582] = 32'hFFFFFFF0;
    // rom_array[1583] = 32'hFFFFFFF0;
    // rom_array[1584] = 32'h00000f99;
    // rom_array[1585] = 32'hFFFFFFF0;
    // rom_array[1586] = 32'h00000fa1;
    // rom_array[1587] = 32'hFFFFFFF0;
    // rom_array[1588] = 32'h00000fa9;
    // rom_array[1589] = 32'hFFFFFFF0;
    // rom_array[1590] = 32'h00000fb1;
    // rom_array[1591] = 32'hFFFFFFF0;
    // rom_array[1592] = 32'h00000fb9;
    // rom_array[1593] = 32'hFFFFFFF0;
    // rom_array[1594] = 32'hFFFFFFF0;
    // rom_array[1595] = 32'hFFFFFFF0;
    // rom_array[1596] = 32'h00000fc1;
    // rom_array[1597] = 32'hFFFFFFF0;
    // rom_array[1598] = 32'hFFFFFFF0;
    // rom_array[1599] = 32'hFFFFFFF0;
    // rom_array[1600] = 32'hFFFFFFF0;
    // rom_array[1601] = 32'hFFFFFFF0;
    // rom_array[1602] = 32'h00000fc9;
    // rom_array[1603] = 32'hFFFFFFF0;
    // rom_array[1604] = 32'h00000fd1;
    // rom_array[1605] = 32'hFFFFFFF0;
    // rom_array[1606] = 32'hFFFFFFF0;
    // rom_array[1607] = 32'hFFFFFFF0;
    // rom_array[1608] = 32'hFFFFFFF0;
    // rom_array[1609] = 32'hFFFFFFF0;
    // rom_array[1610] = 32'hFFFFFFF0;
    // rom_array[1611] = 32'hFFFFFFF0;
    // rom_array[1612] = 32'h00000fd9;
    // rom_array[1613] = 32'hFFFFFFF0;
    // rom_array[1614] = 32'hFFFFFFF0;
    // rom_array[1615] = 32'hFFFFFFF0;
    // rom_array[1616] = 32'h00000fe1;
    // rom_array[1617] = 32'hFFFFFFF0;
    // rom_array[1618] = 32'h00000fe9;
    // rom_array[1619] = 32'hFFFFFFF0;
    // rom_array[1620] = 32'hFFFFFFF0;
    // rom_array[1621] = 32'hFFFFFFF0;
    // rom_array[1622] = 32'h00000ff1;
    // rom_array[1623] = 32'hFFFFFFF0;
    // rom_array[1624] = 32'h00000ff9;
    // rom_array[1625] = 32'hFFFFFFF0;
    // rom_array[1626] = 32'hFFFFFFF0;
    // rom_array[1627] = 32'hFFFFFFF0;
    // rom_array[1628] = 32'h00001001;
    // rom_array[1629] = 32'hFFFFFFF0;
    // rom_array[1630] = 32'hFFFFFFF0;
    // rom_array[1631] = 32'hFFFFFFF0;
    // rom_array[1632] = 32'h00001009;
    // rom_array[1633] = 32'hFFFFFFF0;
    // rom_array[1634] = 32'h00001011;
    // rom_array[1635] = 32'hFFFFFFF0;
    // rom_array[1636] = 32'h00001019;
    // rom_array[1637] = 32'hFFFFFFF0;
    // rom_array[1638] = 32'h00001021;
    // rom_array[1639] = 32'hFFFFFFF0;
    // rom_array[1640] = 32'hFFFFFFF0;
    // rom_array[1641] = 32'hFFFFFFF0;
    // rom_array[1642] = 32'hFFFFFFF0;
    // rom_array[1643] = 32'hFFFFFFF0;
    // rom_array[1644] = 32'h00001029;
    // rom_array[1645] = 32'hFFFFFFF0;
    // rom_array[1646] = 32'hFFFFFFF0;
    // rom_array[1647] = 32'hFFFFFFF0;
    // rom_array[1648] = 32'h00001031;
    // rom_array[1649] = 32'hFFFFFFF0;
    // rom_array[1650] = 32'h00001039;
    // rom_array[1651] = 32'hFFFFFFF0;
    // rom_array[1652] = 32'h00001041;
    // rom_array[1653] = 32'hFFFFFFF0;
    // rom_array[1654] = 32'h00001049;
    // rom_array[1655] = 32'hFFFFFFF0;
    // rom_array[1656] = 32'h00001051;
    // rom_array[1657] = 32'hFFFFFFF0;
    // rom_array[1658] = 32'hFFFFFFF0;
    // rom_array[1659] = 32'hFFFFFFF0;
    // rom_array[1660] = 32'h00001059;
    // rom_array[1661] = 32'hFFFFFFF0;
    // rom_array[1662] = 32'hFFFFFFF0;
    // rom_array[1663] = 32'hFFFFFFF0;
    // rom_array[1664] = 32'h00001061;
    // rom_array[1665] = 32'hFFFFFFF0;
    // rom_array[1666] = 32'h00001069;
    // rom_array[1667] = 32'hFFFFFFF0;
    // rom_array[1668] = 32'h00001071;
    // rom_array[1669] = 32'hFFFFFFF0;
    // rom_array[1670] = 32'h00001079;
    // rom_array[1671] = 32'hFFFFFFF0;
    // rom_array[1672] = 32'h00001081;
    // rom_array[1673] = 32'hFFFFFFF0;
    // rom_array[1674] = 32'hFFFFFFF0;
    // rom_array[1675] = 32'hFFFFFFF0;
    // rom_array[1676] = 32'h00001089;
    // rom_array[1677] = 32'hFFFFFFF0;
    // rom_array[1678] = 32'hFFFFFFF0;
    // rom_array[1679] = 32'hFFFFFFF0;
    // rom_array[1680] = 32'h00001091;
    // rom_array[1681] = 32'hFFFFFFF0;
    // rom_array[1682] = 32'h00001099;
    // rom_array[1683] = 32'hFFFFFFF0;
    // rom_array[1684] = 32'h000010a1;
    // rom_array[1685] = 32'hFFFFFFF0;
    // rom_array[1686] = 32'h000010a9;
    // rom_array[1687] = 32'hFFFFFFF0;
    // rom_array[1688] = 32'h000010b1;
    // rom_array[1689] = 32'hFFFFFFF0;
    // rom_array[1690] = 32'hFFFFFFF0;
    // rom_array[1691] = 32'hFFFFFFF0;
    // rom_array[1692] = 32'hFFFFFFF0;
    // rom_array[1693] = 32'hFFFFFFF0;
    // rom_array[1694] = 32'hFFFFFFF0;
    // rom_array[1695] = 32'hFFFFFFF0;
    // rom_array[1696] = 32'h000010b9;
    // rom_array[1697] = 32'hFFFFFFF0;
    // rom_array[1698] = 32'hFFFFFFF0;
    // rom_array[1699] = 32'hFFFFFFF0;
    // rom_array[1700] = 32'hFFFFFFF0;
    // rom_array[1701] = 32'hFFFFFFF0;
    // rom_array[1702] = 32'h000010c1;
    // rom_array[1703] = 32'hFFFFFFF0;
    // rom_array[1704] = 32'h000010c9;
    // rom_array[1705] = 32'hFFFFFFF0;
    // rom_array[1706] = 32'hFFFFFFF0;
    // rom_array[1707] = 32'hFFFFFFF0;
    // rom_array[1708] = 32'h000010d1;
    // rom_array[1709] = 32'hFFFFFFF0;
    // rom_array[1710] = 32'hFFFFFFF0;
    // rom_array[1711] = 32'hFFFFFFF0;
    // rom_array[1712] = 32'h000010d9;
    // rom_array[1713] = 32'hFFFFFFF0;
    // rom_array[1714] = 32'h000010e1;
    // rom_array[1715] = 32'hFFFFFFF0;
    // rom_array[1716] = 32'h000010e9;
    // rom_array[1717] = 32'hFFFFFFF0;
    // rom_array[1718] = 32'h000010f1;
    // rom_array[1719] = 32'hFFFFFFF0;
    // rom_array[1720] = 32'hFFFFFFF0;
    // rom_array[1721] = 32'hFFFFFFF0;
    // rom_array[1722] = 32'hFFFFFFF0;
    // rom_array[1723] = 32'hFFFFFFF0;
    // rom_array[1724] = 32'h000010f9;
    // rom_array[1725] = 32'hFFFFFFF0;
    // rom_array[1726] = 32'hFFFFFFF0;
    // rom_array[1727] = 32'hFFFFFFF0;
    // rom_array[1728] = 32'hFFFFFFF0;
    // rom_array[1729] = 32'hFFFFFFF0;
    // rom_array[1730] = 32'h00001101;
    // rom_array[1731] = 32'hFFFFFFF0;
    // rom_array[1732] = 32'hFFFFFFF0;
    // rom_array[1733] = 32'hFFFFFFF0;
    // rom_array[1734] = 32'hFFFFFFF0;
    // rom_array[1735] = 32'hFFFFFFF0;
    // rom_array[1736] = 32'hFFFFFFF0;
    // rom_array[1737] = 32'hFFFFFFF0;
    // rom_array[1738] = 32'hFFFFFFF0;
    // rom_array[1739] = 32'h00001109;
    // rom_array[1740] = 32'hFFFFFFF0;
    // rom_array[1741] = 32'hFFFFFFF0;
    // rom_array[1742] = 32'hFFFFFFF0;
    // rom_array[1743] = 32'hFFFFFFF0;
    // rom_array[1744] = 32'hFFFFFFF0;
    // rom_array[1745] = 32'h00001111;
    // rom_array[1746] = 32'hFFFFFFF0;
    // rom_array[1747] = 32'h00001119;
    // rom_array[1748] = 32'hFFFFFFF0;
    // rom_array[1749] = 32'hFFFFFFF0;
    // rom_array[1750] = 32'hFFFFFFF0;
    // rom_array[1751] = 32'hFFFFFFF0;
    // rom_array[1752] = 32'hFFFFFFF0;
    // rom_array[1753] = 32'hFFFFFFF0;
    // rom_array[1754] = 32'hFFFFFFF0;
    // rom_array[1755] = 32'h00001121;
    // rom_array[1756] = 32'hFFFFFFF0;
    // rom_array[1757] = 32'hFFFFFFF0;
    // rom_array[1758] = 32'hFFFFFFF0;
    // rom_array[1759] = 32'h00001129;
    // rom_array[1760] = 32'hFFFFFFF0;
    // rom_array[1761] = 32'h00001131;
    // rom_array[1762] = 32'hFFFFFFF0;
    // rom_array[1763] = 32'h00001139;
    // rom_array[1764] = 32'hFFFFFFF0;
    // rom_array[1765] = 32'h00001141;
    // rom_array[1766] = 32'hFFFFFFF0;
    // rom_array[1767] = 32'h00001149;
    // rom_array[1768] = 32'hFFFFFFF0;
    // rom_array[1769] = 32'hFFFFFFF0;
    // rom_array[1770] = 32'hFFFFFFF0;
    // rom_array[1771] = 32'h00001151;
    // rom_array[1772] = 32'hFFFFFFF0;
    // rom_array[1773] = 32'hFFFFFFF0;
    // rom_array[1774] = 32'hFFFFFFF0;
    // rom_array[1775] = 32'h00001159;
    // rom_array[1776] = 32'hFFFFFFF0;
    // rom_array[1777] = 32'h00001161;
    // rom_array[1778] = 32'hFFFFFFF0;
    // rom_array[1779] = 32'h00001169;
    // rom_array[1780] = 32'hFFFFFFF0;
    // rom_array[1781] = 32'h00001171;
    // rom_array[1782] = 32'hFFFFFFF0;
    // rom_array[1783] = 32'h00001179;
    // rom_array[1784] = 32'hFFFFFFF0;
    // rom_array[1785] = 32'hFFFFFFF0;
    // rom_array[1786] = 32'hFFFFFFF0;
    // rom_array[1787] = 32'h00001181;
    // rom_array[1788] = 32'hFFFFFFF0;
    // rom_array[1789] = 32'hFFFFFFF0;
    // rom_array[1790] = 32'hFFFFFFF0;
    // rom_array[1791] = 32'hFFFFFFF0;
    // rom_array[1792] = 32'hFFFFFFF0;
    // rom_array[1793] = 32'h00001189;
    // rom_array[1794] = 32'hFFFFFFF0;
    // rom_array[1795] = 32'h00001191;
    // rom_array[1796] = 32'hFFFFFFF0;
    // rom_array[1797] = 32'hFFFFFFF0;
    // rom_array[1798] = 32'hFFFFFFF0;
    // rom_array[1799] = 32'hFFFFFFF0;
    // rom_array[1800] = 32'hFFFFFFF0;
    // rom_array[1801] = 32'hFFFFFFF0;
    // rom_array[1802] = 32'hFFFFFFF0;
    // rom_array[1803] = 32'h00001199;
    // rom_array[1804] = 32'hFFFFFFF0;
    // rom_array[1805] = 32'hFFFFFFF0;
    // rom_array[1806] = 32'hFFFFFFF0;
    // rom_array[1807] = 32'h000011a1;
    // rom_array[1808] = 32'hFFFFFFF0;
    // rom_array[1809] = 32'h000011a9;
    // rom_array[1810] = 32'hFFFFFFF0;
    // rom_array[1811] = 32'hFFFFFFF0;
    // rom_array[1812] = 32'hFFFFFFF0;
    // rom_array[1813] = 32'h000011b1;
    // rom_array[1814] = 32'hFFFFFFF0;
    // rom_array[1815] = 32'h000011b9;
    // rom_array[1816] = 32'hFFFFFFF0;
    // rom_array[1817] = 32'hFFFFFFF0;
    // rom_array[1818] = 32'hFFFFFFF0;
    // rom_array[1819] = 32'h000011c1;
    // rom_array[1820] = 32'hFFFFFFF0;
    // rom_array[1821] = 32'hFFFFFFF0;
    // rom_array[1822] = 32'hFFFFFFF0;
    // rom_array[1823] = 32'h000011c9;
    // rom_array[1824] = 32'hFFFFFFF0;
    // rom_array[1825] = 32'h000011d1;
    // rom_array[1826] = 32'hFFFFFFF0;
    // rom_array[1827] = 32'h000011d9;
    // rom_array[1828] = 32'hFFFFFFF0;
    // rom_array[1829] = 32'h000011e1;
    // rom_array[1830] = 32'hFFFFFFF0;
    // rom_array[1831] = 32'hFFFFFFF0;
    // rom_array[1832] = 32'hFFFFFFF0;
    // rom_array[1833] = 32'hFFFFFFF0;
    // rom_array[1834] = 32'hFFFFFFF0;
    // rom_array[1835] = 32'h000011e9;
    // rom_array[1836] = 32'hFFFFFFF0;
    // rom_array[1837] = 32'hFFFFFFF0;
    // rom_array[1838] = 32'hFFFFFFF0;
    // rom_array[1839] = 32'h000011f1;
    // rom_array[1840] = 32'hFFFFFFF0;
    // rom_array[1841] = 32'h000011f9;
    // rom_array[1842] = 32'hFFFFFFF0;
    // rom_array[1843] = 32'h00001201;
    // rom_array[1844] = 32'hFFFFFFF0;
    // rom_array[1845] = 32'h00001209;
    // rom_array[1846] = 32'hFFFFFFF0;
    // rom_array[1847] = 32'h00001211;
    // rom_array[1848] = 32'hFFFFFFF0;
    // rom_array[1849] = 32'hFFFFFFF0;
    // rom_array[1850] = 32'hFFFFFFF0;
    // rom_array[1851] = 32'h00001219;
    // rom_array[1852] = 32'hFFFFFFF0;
    // rom_array[1853] = 32'hFFFFFFF0;
    // rom_array[1854] = 32'hFFFFFFF0;
    // rom_array[1855] = 32'h00001221;
    // rom_array[1856] = 32'hFFFFFFF0;
    // rom_array[1857] = 32'h00001229;
    // rom_array[1858] = 32'hFFFFFFF0;
    // rom_array[1859] = 32'h00001231;
    // rom_array[1860] = 32'hFFFFFFF0;
    // rom_array[1861] = 32'h00001239;
    // rom_array[1862] = 32'hFFFFFFF0;
    // rom_array[1863] = 32'h00001241;
    // rom_array[1864] = 32'hFFFFFFF0;
    // rom_array[1865] = 32'hFFFFFFF0;
    // rom_array[1866] = 32'hFFFFFFF0;
    // rom_array[1867] = 32'h00001249;
    // rom_array[1868] = 32'hFFFFFFF0;
    // rom_array[1869] = 32'hFFFFFFF0;
    // rom_array[1870] = 32'hFFFFFFF0;
    // rom_array[1871] = 32'h00001251;
    // rom_array[1872] = 32'hFFFFFFF0;
    // rom_array[1873] = 32'h00001259;
    // rom_array[1874] = 32'hFFFFFFF0;
    // rom_array[1875] = 32'h00001261;
    // rom_array[1876] = 32'hFFFFFFF0;
    // rom_array[1877] = 32'h00001269;
    // rom_array[1878] = 32'hFFFFFFF0;
    // rom_array[1879] = 32'h00001271;
    // rom_array[1880] = 32'hFFFFFFF0;
    // rom_array[1881] = 32'hFFFFFFF0;
    // rom_array[1882] = 32'hFFFFFFF0;
    // rom_array[1883] = 32'hFFFFFFF0;
    // rom_array[1884] = 32'hFFFFFFF0;
    // rom_array[1885] = 32'hFFFFFFF0;
    // rom_array[1886] = 32'hFFFFFFF0;
    // rom_array[1887] = 32'h00001279;
    // rom_array[1888] = 32'hFFFFFFF0;
    // rom_array[1889] = 32'hFFFFFFF0;
    // rom_array[1890] = 32'hFFFFFFF0;
    // rom_array[1891] = 32'hFFFFFFF0;
    // rom_array[1892] = 32'hFFFFFFF0;
    // rom_array[1893] = 32'h00001281;
    // rom_array[1894] = 32'hFFFFFFF0;
    // rom_array[1895] = 32'h00001289;
    // rom_array[1896] = 32'hFFFFFFF0;
    // rom_array[1897] = 32'hFFFFFFF0;
    // rom_array[1898] = 32'hFFFFFFF0;
    // rom_array[1899] = 32'h00001291;
    // rom_array[1900] = 32'hFFFFFFF0;
    // rom_array[1901] = 32'hFFFFFFF0;
    // rom_array[1902] = 32'hFFFFFFF0;
    // rom_array[1903] = 32'h00001299;
    // rom_array[1904] = 32'hFFFFFFF0;
    // rom_array[1905] = 32'h000012a1;
    // rom_array[1906] = 32'hFFFFFFF0;
    // rom_array[1907] = 32'h000012a9;
    // rom_array[1908] = 32'hFFFFFFF0;
    // rom_array[1909] = 32'h000012b1;
    // rom_array[1910] = 32'hFFFFFFF0;
    // rom_array[1911] = 32'hFFFFFFF0;
    // rom_array[1912] = 32'hFFFFFFF0;
    // rom_array[1913] = 32'hFFFFFFF0;
    // rom_array[1914] = 32'hFFFFFFF0;
    // rom_array[1915] = 32'h000012b9;
    // rom_array[1916] = 32'hFFFFFFF0;
    // rom_array[1917] = 32'hFFFFFFF0;
    // rom_array[1918] = 32'hFFFFFFF0;
    // rom_array[1919] = 32'hFFFFFFF0;
    // rom_array[1920] = 32'hFFFFFFF0;
    // rom_array[1921] = 32'h000012c1;
    // rom_array[1922] = 32'hFFFFFFF0;
    // rom_array[1923] = 32'hFFFFFFF0;
    // rom_array[1924] = 32'hFFFFFFF0;
    // rom_array[1925] = 32'hFFFFFFF0;
    // rom_array[1926] = 32'hFFFFFFF0;
    // rom_array[1927] = 32'hFFFFFFF0;
    // rom_array[1928] = 32'hFFFFFFF0;
    // rom_array[1929] = 32'hFFFFFFF0;
    // rom_array[1930] = 32'h000012c9;
    // rom_array[1931] = 32'hFFFFFFF0;
    // rom_array[1932] = 32'h000012d1;
    // rom_array[1933] = 32'hFFFFFFF0;
    // rom_array[1934] = 32'hFFFFFFF0;
    // rom_array[1935] = 32'hFFFFFFF0;
    // rom_array[1936] = 32'hFFFFFFF0;
    // rom_array[1937] = 32'hFFFFFFF0;
    // rom_array[1938] = 32'h000012d9;
    // rom_array[1939] = 32'hFFFFFFF0;
    // rom_array[1940] = 32'hFFFFFFF0;
    // rom_array[1941] = 32'hFFFFFFF0;
    // rom_array[1942] = 32'hFFFFFFF0;
    // rom_array[1943] = 32'hFFFFFFF0;
    // rom_array[1944] = 32'hFFFFFFF0;
    // rom_array[1945] = 32'hFFFFFFF0;
    // rom_array[1946] = 32'h000012e1;
    // rom_array[1947] = 32'hFFFFFFF0;
    // rom_array[1948] = 32'h000012e9;
    // rom_array[1949] = 32'hFFFFFFF0;
    // rom_array[1950] = 32'h000012f1;
    // rom_array[1951] = 32'hFFFFFFF0;
    // rom_array[1952] = 32'h000012f9;
    // rom_array[1953] = 32'hFFFFFFF0;
    // rom_array[1954] = 32'h00001301;
    // rom_array[1955] = 32'hFFFFFFF0;
    // rom_array[1956] = 32'hFFFFFFF0;
    // rom_array[1957] = 32'hFFFFFFF0;
    // rom_array[1958] = 32'h00001309;
    // rom_array[1959] = 32'hFFFFFFF0;
    // rom_array[1960] = 32'hFFFFFFF0;
    // rom_array[1961] = 32'hFFFFFFF0;
    // rom_array[1962] = 32'h00001311;
    // rom_array[1963] = 32'hFFFFFFF0;
    // rom_array[1964] = 32'h00001319;
    // rom_array[1965] = 32'hFFFFFFF0;
    // rom_array[1966] = 32'h00001321;
    // rom_array[1967] = 32'hFFFFFFF0;
    // rom_array[1968] = 32'h00001329;
    // rom_array[1969] = 32'hFFFFFFF0;
    // rom_array[1970] = 32'h00001331;
    // rom_array[1971] = 32'hFFFFFFF0;
    // rom_array[1972] = 32'hFFFFFFF0;
    // rom_array[1973] = 32'hFFFFFFF0;
    // rom_array[1974] = 32'h00001339;
    // rom_array[1975] = 32'hFFFFFFF0;
    // rom_array[1976] = 32'hFFFFFFF0;
    // rom_array[1977] = 32'hFFFFFFF0;
    // rom_array[1978] = 32'h00001341;
    // rom_array[1979] = 32'hFFFFFFF0;
    // rom_array[1980] = 32'h00001349;
    // rom_array[1981] = 32'hFFFFFFF0;
    // rom_array[1982] = 32'hFFFFFFF0;
    // rom_array[1983] = 32'hFFFFFFF0;
    // rom_array[1984] = 32'hFFFFFFF0;
    // rom_array[1985] = 32'hFFFFFFF0;
    // rom_array[1986] = 32'hFFFFFFF0;
    // rom_array[1987] = 32'hFFFFFFF0;
    // rom_array[1988] = 32'h00001351;
    // rom_array[1989] = 32'hFFFFFFF0;
    // rom_array[1990] = 32'h00001359;
    // rom_array[1991] = 32'hFFFFFFF0;
    // rom_array[1992] = 32'h00001361;
    // rom_array[1993] = 32'hFFFFFFF0;
    // rom_array[1994] = 32'h00001369;
    // rom_array[1995] = 32'hFFFFFFF0;
    // rom_array[1996] = 32'hFFFFFFF0;
    // rom_array[1997] = 32'hFFFFFFF0;
    // rom_array[1998] = 32'h00001371;
    // rom_array[1999] = 32'hFFFFFFF0;
    // rom_array[2000] = 32'hFFFFFFF0;
    // rom_array[2001] = 32'hFFFFFFF0;
    // rom_array[2002] = 32'h00001379;
    // rom_array[2003] = 32'hFFFFFFF0;
    // rom_array[2004] = 32'h00001381;
    // rom_array[2005] = 32'hFFFFFFF0;
    // rom_array[2006] = 32'hFFFFFFF0;
    // rom_array[2007] = 32'hFFFFFFF0;
    // rom_array[2008] = 32'h00001389;
    // rom_array[2009] = 32'hFFFFFFF0;
    // rom_array[2010] = 32'h00001391;
    // rom_array[2011] = 32'hFFFFFFF0;
    // rom_array[2012] = 32'hFFFFFFF0;
    // rom_array[2013] = 32'hFFFFFFF0;
    // rom_array[2014] = 32'h00001399;
    // rom_array[2015] = 32'hFFFFFFF0;
    // rom_array[2016] = 32'hFFFFFFF0;
    // rom_array[2017] = 32'hFFFFFFF0;
    // rom_array[2018] = 32'h000013a1;
    // rom_array[2019] = 32'hFFFFFFF0;
    // rom_array[2020] = 32'h000013a9;
    // rom_array[2021] = 32'hFFFFFFF0;
    // rom_array[2022] = 32'h000013b1;
    // rom_array[2023] = 32'hFFFFFFF0;
    // rom_array[2024] = 32'h000013b9;
    // rom_array[2025] = 32'hFFFFFFF0;
    // rom_array[2026] = 32'h000013c1;
    // rom_array[2027] = 32'hFFFFFFF0;
    // rom_array[2028] = 32'hFFFFFFF0;
    // rom_array[2029] = 32'hFFFFFFF0;
    // rom_array[2030] = 32'h000013c9;
    // rom_array[2031] = 32'hFFFFFFF0;
    // rom_array[2032] = 32'hFFFFFFF0;
    // rom_array[2033] = 32'hFFFFFFF0;
    // rom_array[2034] = 32'h000013d1;
    // rom_array[2035] = 32'hFFFFFFF0;
    // rom_array[2036] = 32'h000013d9;
    // rom_array[2037] = 32'hFFFFFFF0;
    // rom_array[2038] = 32'h000013e1;
    // rom_array[2039] = 32'hFFFFFFF0;
    // rom_array[2040] = 32'h000013e9;
    // rom_array[2041] = 32'hFFFFFFF0;
    // rom_array[2042] = 32'h000013f1;
    // rom_array[2043] = 32'hFFFFFFF0;
    // rom_array[2044] = 32'hFFFFFFF0;
    // rom_array[2045] = 32'hFFFFFFF0;
    // rom_array[2046] = 32'h000013f9;
    // rom_array[2047] = 32'hFFFFFFF0;
    // rom_array[2048] = 32'hFFFFFFF0;
    // rom_array[2049] = 32'hFFFFFFF0;
    // rom_array[2050] = 32'h00001401;
    // rom_array[2051] = 32'hFFFFFFF0;
    // rom_array[2052] = 32'h00001409;
    // rom_array[2053] = 32'hFFFFFFF0;
    // rom_array[2054] = 32'h00001411;
    // rom_array[2055] = 32'hFFFFFFF0;
    // rom_array[2056] = 32'h00001419;
    // rom_array[2057] = 32'hFFFFFFF0;
    // rom_array[2058] = 32'h00001421;
    // rom_array[2059] = 32'hFFFFFFF0;
    // rom_array[2060] = 32'hFFFFFFF0;
    // rom_array[2061] = 32'hFFFFFFF0;
    // rom_array[2062] = 32'h00001429;
    // rom_array[2063] = 32'hFFFFFFF0;
    // rom_array[2064] = 32'hFFFFFFF0;
    // rom_array[2065] = 32'hFFFFFFF0;
    // rom_array[2066] = 32'hFFFFFFF0;
    // rom_array[2067] = 32'hFFFFFFF0;
    // rom_array[2068] = 32'hFFFFFFF0;
    // rom_array[2069] = 32'hFFFFFFF0;
    // rom_array[2070] = 32'h00001431;
    // rom_array[2071] = 32'hFFFFFFF0;
    // rom_array[2072] = 32'h00001439;
    // rom_array[2073] = 32'hFFFFFFF0;
    // rom_array[2074] = 32'hFFFFFFF0;
    // rom_array[2075] = 32'hFFFFFFF0;
    // rom_array[2076] = 32'hFFFFFFF0;
    // rom_array[2077] = 32'hFFFFFFF0;
    // rom_array[2078] = 32'h00001441;
    // rom_array[2079] = 32'hFFFFFFF0;
    // rom_array[2080] = 32'hFFFFFFF0;
    // rom_array[2081] = 32'hFFFFFFF0;
    // rom_array[2082] = 32'h00001449;
    // rom_array[2083] = 32'hFFFFFFF0;
    // rom_array[2084] = 32'h00001451;
    // rom_array[2085] = 32'hFFFFFFF0;
    // rom_array[2086] = 32'hFFFFFFF0;
    // rom_array[2087] = 32'hFFFFFFF0;
    // rom_array[2088] = 32'hFFFFFFF0;
    // rom_array[2089] = 32'hFFFFFFF0;
    // rom_array[2090] = 32'h00001459;
    // rom_array[2091] = 32'hFFFFFFF0;
    // rom_array[2092] = 32'hFFFFFFF0;
    // rom_array[2093] = 32'hFFFFFFF0;
    // rom_array[2094] = 32'hFFFFFFF0;
    // rom_array[2095] = 32'hFFFFFFF0;
    // rom_array[2096] = 32'hFFFFFFF0;
    // rom_array[2097] = 32'h00001461;
    // rom_array[2098] = 32'hFFFFFFF0;
    // rom_array[2099] = 32'h00001469;
    // rom_array[2100] = 32'hFFFFFFF0;
    // rom_array[2101] = 32'hFFFFFFF0;
    // rom_array[2102] = 32'hFFFFFFF0;
    // rom_array[2103] = 32'hFFFFFFF0;
    // rom_array[2104] = 32'hFFFFFFF0;
    // rom_array[2105] = 32'h00001471;
    // rom_array[2106] = 32'hFFFFFFF0;
    // rom_array[2107] = 32'hFFFFFFF0;
    // rom_array[2108] = 32'hFFFFFFF0;
    // rom_array[2109] = 32'hFFFFFFF0;
    // rom_array[2110] = 32'hFFFFFFF0;
    // rom_array[2111] = 32'hFFFFFFF0;
    // rom_array[2112] = 32'hFFFFFFF0;
    // rom_array[2113] = 32'h00001479;
    // rom_array[2114] = 32'hFFFFFFF0;
    // rom_array[2115] = 32'h00001481;
    // rom_array[2116] = 32'hFFFFFFF0;
    // rom_array[2117] = 32'h00001489;
    // rom_array[2118] = 32'hFFFFFFF0;
    // rom_array[2119] = 32'h00001491;
    // rom_array[2120] = 32'hFFFFFFF0;
    // rom_array[2121] = 32'h00001499;
    // rom_array[2122] = 32'hFFFFFFF0;
    // rom_array[2123] = 32'hFFFFFFF0;
    // rom_array[2124] = 32'hFFFFFFF0;
    // rom_array[2125] = 32'h000014a1;
    // rom_array[2126] = 32'hFFFFFFF0;
    // rom_array[2127] = 32'hFFFFFFF0;
    // rom_array[2128] = 32'hFFFFFFF0;
    // rom_array[2129] = 32'h000014a9;
    // rom_array[2130] = 32'hFFFFFFF0;
    // rom_array[2131] = 32'h000014b1;
    // rom_array[2132] = 32'hFFFFFFF0;
    // rom_array[2133] = 32'h000014b9;
    // rom_array[2134] = 32'hFFFFFFF0;
    // rom_array[2135] = 32'h000014c1;
    // rom_array[2136] = 32'hFFFFFFF0;
    // rom_array[2137] = 32'h000014c9;
    // rom_array[2138] = 32'hFFFFFFF0;
    // rom_array[2139] = 32'hFFFFFFF0;
    // rom_array[2140] = 32'hFFFFFFF0;
    // rom_array[2141] = 32'h000014d1;
    // rom_array[2142] = 32'hFFFFFFF0;
    // rom_array[2143] = 32'hFFFFFFF0;
    // rom_array[2144] = 32'hFFFFFFF0;
    // rom_array[2145] = 32'h000014d9;
    // rom_array[2146] = 32'hFFFFFFF0;
    // rom_array[2147] = 32'h000014e1;
    // rom_array[2148] = 32'hFFFFFFF0;
    // rom_array[2149] = 32'hFFFFFFF0;
    // rom_array[2150] = 32'hFFFFFFF0;
    // rom_array[2151] = 32'hFFFFFFF0;
    // rom_array[2152] = 32'hFFFFFFF0;
    // rom_array[2153] = 32'hFFFFFFF0;
    // rom_array[2154] = 32'hFFFFFFF0;
    // rom_array[2155] = 32'h000014e9;
    // rom_array[2156] = 32'hFFFFFFF0;
    // rom_array[2157] = 32'h000014f1;
    // rom_array[2158] = 32'hFFFFFFF0;
    // rom_array[2159] = 32'h000014f9;
    // rom_array[2160] = 32'hFFFFFFF0;
    // rom_array[2161] = 32'h00001501;
    // rom_array[2162] = 32'hFFFFFFF0;
    // rom_array[2163] = 32'hFFFFFFF0;
    // rom_array[2164] = 32'hFFFFFFF0;
    // rom_array[2165] = 32'h00001509;
    // rom_array[2166] = 32'hFFFFFFF0;
    // rom_array[2167] = 32'hFFFFFFF0;
    // rom_array[2168] = 32'hFFFFFFF0;
    // rom_array[2169] = 32'h00001511;
    // rom_array[2170] = 32'hFFFFFFF0;
    // rom_array[2171] = 32'h00001519;
    // rom_array[2172] = 32'hFFFFFFF0;
    // rom_array[2173] = 32'hFFFFFFF0;
    // rom_array[2174] = 32'hFFFFFFF0;
    // rom_array[2175] = 32'h00001521;
    // rom_array[2176] = 32'hFFFFFFF0;
    // rom_array[2177] = 32'h00001529;
    // rom_array[2178] = 32'hFFFFFFF0;
    // rom_array[2179] = 32'hFFFFFFF0;
    // rom_array[2180] = 32'hFFFFFFF0;
    // rom_array[2181] = 32'h00001531;
    // rom_array[2182] = 32'hFFFFFFF0;
    // rom_array[2183] = 32'hFFFFFFF0;
    // rom_array[2184] = 32'hFFFFFFF0;
    // rom_array[2185] = 32'h00001539;
    // rom_array[2186] = 32'hFFFFFFF0;
    // rom_array[2187] = 32'h00001541;
    // rom_array[2188] = 32'hFFFFFFF0;
    // rom_array[2189] = 32'h00001549;
    // rom_array[2190] = 32'hFFFFFFF0;
    // rom_array[2191] = 32'h00001551;
    // rom_array[2192] = 32'hFFFFFFF0;
    // rom_array[2193] = 32'h00001559;
    // rom_array[2194] = 32'hFFFFFFF0;
    // rom_array[2195] = 32'hFFFFFFF0;
    // rom_array[2196] = 32'hFFFFFFF0;
    // rom_array[2197] = 32'h00001561;
    // rom_array[2198] = 32'hFFFFFFF0;
    // rom_array[2199] = 32'hFFFFFFF0;
    // rom_array[2200] = 32'hFFFFFFF0;
    // rom_array[2201] = 32'h00001569;
    // rom_array[2202] = 32'hFFFFFFF0;
    // rom_array[2203] = 32'h00001571;
    // rom_array[2204] = 32'hFFFFFFF0;
    // rom_array[2205] = 32'h00001579;
    // rom_array[2206] = 32'hFFFFFFF0;
    // rom_array[2207] = 32'h00001581;
    // rom_array[2208] = 32'hFFFFFFF0;
    // rom_array[2209] = 32'h00001589;
    // rom_array[2210] = 32'hFFFFFFF0;
    // rom_array[2211] = 32'hFFFFFFF0;
    // rom_array[2212] = 32'hFFFFFFF0;
    // rom_array[2213] = 32'h00001591;
    // rom_array[2214] = 32'hFFFFFFF0;
    // rom_array[2215] = 32'hFFFFFFF0;
    // rom_array[2216] = 32'hFFFFFFF0;
    // rom_array[2217] = 32'h00001599;
    // rom_array[2218] = 32'hFFFFFFF0;
    // rom_array[2219] = 32'h000015a1;
    // rom_array[2220] = 32'hFFFFFFF0;
    // rom_array[2221] = 32'h000015a9;
    // rom_array[2222] = 32'hFFFFFFF0;
    // rom_array[2223] = 32'h000015b1;
    // rom_array[2224] = 32'hFFFFFFF0;
    // rom_array[2225] = 32'h000015b9;
    // rom_array[2226] = 32'hFFFFFFF0;
    // rom_array[2227] = 32'hFFFFFFF0;
    // rom_array[2228] = 32'hFFFFFFF0;
    // rom_array[2229] = 32'h000015c1;
    // rom_array[2230] = 32'hFFFFFFF0;
    // rom_array[2231] = 32'hFFFFFFF0;
    // rom_array[2232] = 32'hFFFFFFF0;
    // rom_array[2233] = 32'hFFFFFFF0;
    // rom_array[2234] = 32'hFFFFFFF0;
    // rom_array[2235] = 32'hFFFFFFF0;
    // rom_array[2236] = 32'hFFFFFFF0;
    // rom_array[2237] = 32'h000015c9;
    // rom_array[2238] = 32'hFFFFFFF0;
    // rom_array[2239] = 32'h000015d1;
    // rom_array[2240] = 32'hFFFFFFF0;
    // rom_array[2241] = 32'hFFFFFFF0;
    // rom_array[2242] = 32'hFFFFFFF0;
    // rom_array[2243] = 32'hFFFFFFF0;
    // rom_array[2244] = 32'hFFFFFFF0;
    // rom_array[2245] = 32'h000015d9;
    // rom_array[2246] = 32'hFFFFFFF0;
    // rom_array[2247] = 32'hFFFFFFF0;
    // rom_array[2248] = 32'hFFFFFFF0;
    // rom_array[2249] = 32'h000015e1;
    // rom_array[2250] = 32'hFFFFFFF0;
    // rom_array[2251] = 32'h000015e9;
    // rom_array[2252] = 32'hFFFFFFF0;
    // rom_array[2253] = 32'hFFFFFFF0;
    // rom_array[2254] = 32'hFFFFFFF0;
    // rom_array[2255] = 32'hFFFFFFF0;
    // rom_array[2256] = 32'hFFFFFFF0;
    // rom_array[2257] = 32'h000015f1;
    // rom_array[2258] = 32'hFFFFFFF0;
    // rom_array[2259] = 32'hFFFFFFF0;
    // rom_array[2260] = 32'hFFFFFFF0;
    // rom_array[2261] = 32'hFFFFFFF0;
    // rom_array[2262] = 32'hFFFFFFF0;
    // rom_array[2263] = 32'hFFFFFFF0;
    // rom_array[2264] = 32'hFFFFFFF0;
    // rom_array[2265] = 32'hFFFFFFF0;
    // rom_array[2266] = 32'h000015f9;
    // rom_array[2267] = 32'hFFFFFFF0;
    // rom_array[2268] = 32'h00001601;
    // rom_array[2269] = 32'hFFFFFFF0;
    // rom_array[2270] = 32'h00001609;
    // rom_array[2271] = 32'hFFFFFFF0;
    // rom_array[2272] = 32'hFFFFFFF1;
    // rom_array[2273] = 32'hFFFFFFF0;
    // rom_array[2274] = 32'h00001611;
    // rom_array[2275] = 32'hFFFFFFF0;
    // rom_array[2276] = 32'hFFFFFFF0;
    // rom_array[2277] = 32'hFFFFFFF0;
    // rom_array[2278] = 32'h00001619;
    // rom_array[2279] = 32'hFFFFFFF0;
    // rom_array[2280] = 32'hFFFFFFF0;
    // rom_array[2281] = 32'hFFFFFFF0;
    // rom_array[2282] = 32'h00001621;
    // rom_array[2283] = 32'hFFFFFFF0;
    // rom_array[2284] = 32'hFFFFFFF1;
    // rom_array[2285] = 32'hFFFFFFF0;
    // rom_array[2286] = 32'h00001629;
    // rom_array[2287] = 32'hFFFFFFF0;
    // rom_array[2288] = 32'hFFFFFFF1;
    // rom_array[2289] = 32'hFFFFFFF0;
    // rom_array[2290] = 32'h00001631;
    // rom_array[2291] = 32'hFFFFFFF0;
    // rom_array[2292] = 32'hFFFFFFF1;
    // rom_array[2293] = 32'hFFFFFFF0;
    // rom_array[2294] = 32'h00001639;
    // rom_array[2295] = 32'hFFFFFFF0;
    // rom_array[2296] = 32'hFFFFFFF1;
    // rom_array[2297] = 32'hFFFFFFF0;
    // rom_array[2298] = 32'h00001641;
    // rom_array[2299] = 32'hFFFFFFF0;
    // rom_array[2300] = 32'hFFFFFFF0;
    // rom_array[2301] = 32'hFFFFFFF0;
    // rom_array[2302] = 32'h00001649;
    // rom_array[2303] = 32'hFFFFFFF0;
    // rom_array[2304] = 32'h00001651;
    // rom_array[2305] = 32'hFFFFFFF0;
    // rom_array[2306] = 32'hFFFFFFF0;
    // rom_array[2307] = 32'hFFFFFFF0;
    // rom_array[2308] = 32'hFFFFFFF0;
    // rom_array[2309] = 32'hFFFFFFF0;
    // rom_array[2310] = 32'h00001659;
    // rom_array[2311] = 32'hFFFFFFF0;
    // rom_array[2312] = 32'h00001661;
    // rom_array[2313] = 32'hFFFFFFF0;
    // rom_array[2314] = 32'h00001669;
    // rom_array[2315] = 32'hFFFFFFF0;
    // rom_array[2316] = 32'hFFFFFFF1;
    // rom_array[2317] = 32'hFFFFFFF0;
    // rom_array[2318] = 32'h00001671;
    // rom_array[2319] = 32'hFFFFFFF0;
    // rom_array[2320] = 32'h00001679;
    // rom_array[2321] = 32'hFFFFFFF0;
    // rom_array[2322] = 32'hFFFFFFF1;
    // rom_array[2323] = 32'hFFFFFFF0;
    // rom_array[2324] = 32'hFFFFFFF1;
    // rom_array[2325] = 32'hFFFFFFF0;
    // rom_array[2326] = 32'h00001681;
    // rom_array[2327] = 32'hFFFFFFF0;
    // rom_array[2328] = 32'h00001689;
    // rom_array[2329] = 32'hFFFFFFF0;
    // rom_array[2330] = 32'h00001691;
    // rom_array[2331] = 32'hFFFFFFF0;
    // rom_array[2332] = 32'hFFFFFFF1;
    // rom_array[2333] = 32'hFFFFFFF0;
    // rom_array[2334] = 32'h00001699;
    // rom_array[2335] = 32'hFFFFFFF0;
    // rom_array[2336] = 32'h000016a1;
    // rom_array[2337] = 32'hFFFFFFF0;
    // rom_array[2338] = 32'h000016a9;
    // rom_array[2339] = 32'hFFFFFFF0;
    // rom_array[2340] = 32'hFFFFFFF0;
    // rom_array[2341] = 32'hFFFFFFF0;
    // rom_array[2342] = 32'h000016b1;
    // rom_array[2343] = 32'hFFFFFFF0;
    // rom_array[2344] = 32'hFFFFFFF0;
    // rom_array[2345] = 32'hFFFFFFF0;
    // rom_array[2346] = 32'hFFFFFFF0;
    // rom_array[2347] = 32'hFFFFFFF0;
    // rom_array[2348] = 32'hFFFFFFF0;
    // rom_array[2349] = 32'hFFFFFFF0;
    // rom_array[2350] = 32'h000016b9;
    // rom_array[2351] = 32'hFFFFFFF0;
    // rom_array[2352] = 32'h000016c1;
    // rom_array[2353] = 32'hFFFFFFF0;
    // rom_array[2354] = 32'hFFFFFFF0;
    // rom_array[2355] = 32'hFFFFFFF0;
    // rom_array[2356] = 32'hFFFFFFF0;
    // rom_array[2357] = 32'hFFFFFFF0;
    // rom_array[2358] = 32'h000016c9;
    // rom_array[2359] = 32'hFFFFFFF0;
    // rom_array[2360] = 32'h000016d1;
    // rom_array[2361] = 32'hFFFFFFF0;
    // rom_array[2362] = 32'hFFFFFFF0;
    // rom_array[2363] = 32'hFFFFFFF0;
    // rom_array[2364] = 32'hFFFFFFF0;
    // rom_array[2365] = 32'hFFFFFFF0;
    // rom_array[2366] = 32'h000016d9;
    // rom_array[2367] = 32'hFFFFFFF0;
    // rom_array[2368] = 32'h000016e1;
    // rom_array[2369] = 32'hFFFFFFF0;
    // rom_array[2370] = 32'h000016e9;
    // rom_array[2371] = 32'hFFFFFFF0;
    // rom_array[2372] = 32'hFFFFFFF1;
    // rom_array[2373] = 32'hFFFFFFF0;
    // rom_array[2374] = 32'h000016f1;
    // rom_array[2375] = 32'hFFFFFFF0;
    // rom_array[2376] = 32'h000016f9;
    // rom_array[2377] = 32'hFFFFFFF0;
    // rom_array[2378] = 32'hFFFFFFF1;
    // rom_array[2379] = 32'hFFFFFFF0;
    // rom_array[2380] = 32'h00001701;
    // rom_array[2381] = 32'hFFFFFFF0;
    // rom_array[2382] = 32'h00001709;
    // rom_array[2383] = 32'hFFFFFFF0;
    // rom_array[2384] = 32'h00001711;
    // rom_array[2385] = 32'hFFFFFFF0;
    // rom_array[2386] = 32'hFFFFFFF1;
    // rom_array[2387] = 32'hFFFFFFF0;
    // rom_array[2388] = 32'hFFFFFFF1;
    // rom_array[2389] = 32'hFFFFFFF0;
    // rom_array[2390] = 32'h00001719;
    // rom_array[2391] = 32'hFFFFFFF0;
    // rom_array[2392] = 32'h00001721;
    // rom_array[2393] = 32'hFFFFFFF0;
    // rom_array[2394] = 32'hFFFFFFF0;
    // rom_array[2395] = 32'hFFFFFFF0;
    // rom_array[2396] = 32'h00001729;
    // rom_array[2397] = 32'hFFFFFFF0;
    // rom_array[2398] = 32'hFFFFFFF0;
    // rom_array[2399] = 32'hFFFFFFF0;
    // rom_array[2400] = 32'h00001731;
    // rom_array[2401] = 32'hFFFFFFF0;
    // rom_array[2402] = 32'hFFFFFFF1;
    // rom_array[2403] = 32'hFFFFFFF0;
    // rom_array[2404] = 32'hFFFFFFF1;
    // rom_array[2405] = 32'hFFFFFFF0;
    // rom_array[2406] = 32'h00001739;
    // rom_array[2407] = 32'hFFFFFFF0;
    // rom_array[2408] = 32'h00001741;
    // rom_array[2409] = 32'hFFFFFFF0;
    // rom_array[2410] = 32'hFFFFFFF0;
    // rom_array[2411] = 32'hFFFFFFF0;
    // rom_array[2412] = 32'h00001749;
    // rom_array[2413] = 32'hFFFFFFF0;
    // rom_array[2414] = 32'hFFFFFFF0;
    // rom_array[2415] = 32'hFFFFFFF0;
    // rom_array[2416] = 32'h00001751;
    // rom_array[2417] = 32'hFFFFFFF0;
    // rom_array[2418] = 32'h00001759;
    // rom_array[2419] = 32'hFFFFFFF0;
    // rom_array[2420] = 32'h00001761;
    // rom_array[2421] = 32'hFFFFFFF0;
    // rom_array[2422] = 32'h00001769;
    // rom_array[2423] = 32'hFFFFFFF0;
    // rom_array[2424] = 32'h00001771;
    // rom_array[2425] = 32'hFFFFFFF0;
    // rom_array[2426] = 32'hFFFFFFF0;
    // rom_array[2427] = 32'hFFFFFFF0;
    // rom_array[2428] = 32'h00001779;
    // rom_array[2429] = 32'hFFFFFFF0;
    // rom_array[2430] = 32'hFFFFFFF0;
    // rom_array[2431] = 32'hFFFFFFF0;
    // rom_array[2432] = 32'h00001781;
    // rom_array[2433] = 32'hFFFFFFF0;
    // rom_array[2434] = 32'hFFFFFFF1;
    // rom_array[2435] = 32'hFFFFFFF0;
    // rom_array[2436] = 32'hFFFFFFF1;
    // rom_array[2437] = 32'hFFFFFFF0;
    // rom_array[2438] = 32'hFFFFFFF1;
    // rom_array[2439] = 32'hFFFFFFF0;
    // rom_array[2440] = 32'hFFFFFFF1;
    // rom_array[2441] = 32'hFFFFFFF0;
    // rom_array[2442] = 32'h00001789;
    // rom_array[2443] = 32'hFFFFFFF0;
    // rom_array[2444] = 32'h00001791;
    // rom_array[2445] = 32'hFFFFFFF0;
    // rom_array[2446] = 32'h00001799;
    // rom_array[2447] = 32'hFFFFFFF0;
    // rom_array[2448] = 32'hFFFFFFF1;
    // rom_array[2449] = 32'hFFFFFFF0;
    // rom_array[2450] = 32'h000017a1;
    // rom_array[2451] = 32'hFFFFFFF0;
    // rom_array[2452] = 32'h000017a9;
    // rom_array[2453] = 32'hFFFFFFF0;
    // rom_array[2454] = 32'hFFFFFFF0;
    // rom_array[2455] = 32'hFFFFFFF0;
    // rom_array[2456] = 32'hFFFFFFF0;
    // rom_array[2457] = 32'hFFFFFFF0;
    // rom_array[2458] = 32'h000017b1;
    // rom_array[2459] = 32'hFFFFFFF0;
    // rom_array[2460] = 32'h000017b9;
    // rom_array[2461] = 32'hFFFFFFF0;
    // rom_array[2462] = 32'hFFFFFFF1;
    // rom_array[2463] = 32'hFFFFFFF0;
    // rom_array[2464] = 32'h000017c1;
    // rom_array[2465] = 32'hFFFFFFF0;
    // rom_array[2466] = 32'h000017c9;
    // rom_array[2467] = 32'hFFFFFFF0;
    // rom_array[2468] = 32'h000017d1;
    // rom_array[2469] = 32'hFFFFFFF0;
    // rom_array[2470] = 32'h000017d9;
    // rom_array[2471] = 32'hFFFFFFF0;
    // rom_array[2472] = 32'h000017e1;
    // rom_array[2473] = 32'hFFFFFFF0;
    // rom_array[2474] = 32'h000017e9;
    // rom_array[2475] = 32'hFFFFFFF0;
    // rom_array[2476] = 32'h000017f1;
    // rom_array[2477] = 32'hFFFFFFF0;
    // rom_array[2478] = 32'hFFFFFFF0;
    // rom_array[2479] = 32'hFFFFFFF0;
    // rom_array[2480] = 32'hFFFFFFF0;
    // rom_array[2481] = 32'hFFFFFFF0;
    // rom_array[2482] = 32'h000017f9;
    // rom_array[2483] = 32'hFFFFFFF0;
    // rom_array[2484] = 32'h00001801;
    // rom_array[2485] = 32'hFFFFFFF0;
    // rom_array[2486] = 32'hFFFFFFF0;
    // rom_array[2487] = 32'hFFFFFFF0;
    // rom_array[2488] = 32'hFFFFFFF0;
    // rom_array[2489] = 32'hFFFFFFF0;
    // rom_array[2490] = 32'h00001809;
    // rom_array[2491] = 32'hFFFFFFF0;
    // rom_array[2492] = 32'h00001811;
    // rom_array[2493] = 32'hFFFFFFF0;
    // rom_array[2494] = 32'h00001819;
    // rom_array[2495] = 32'hFFFFFFF0;
    // rom_array[2496] = 32'hFFFFFFF1;
    // rom_array[2497] = 32'hFFFFFFF0;
    // rom_array[2498] = 32'h00001821;
    // rom_array[2499] = 32'hFFFFFFF0;
    // rom_array[2500] = 32'h00001829;
    // rom_array[2501] = 32'hFFFFFFF0;
    // rom_array[2502] = 32'hFFFFFFF0;
    // rom_array[2503] = 32'hFFFFFFF0;
    // rom_array[2504] = 32'hFFFFFFF0;
    // rom_array[2505] = 32'hFFFFFFF0;
    // rom_array[2506] = 32'h00001831;
    // rom_array[2507] = 32'hFFFFFFF0;
    // rom_array[2508] = 32'h00001839;
    // rom_array[2509] = 32'hFFFFFFF0;
    // rom_array[2510] = 32'hFFFFFFF1;
    // rom_array[2511] = 32'hFFFFFFF0;
    // rom_array[2512] = 32'hFFFFFFF1;
    // rom_array[2513] = 32'hFFFFFFF0;
    // rom_array[2514] = 32'h00001841;
    // rom_array[2515] = 32'hFFFFFFF0;
    // rom_array[2516] = 32'h00001849;
    // rom_array[2517] = 32'hFFFFFFF0;
    // rom_array[2518] = 32'hFFFFFFF1;
    // rom_array[2519] = 32'hFFFFFFF0;
    // rom_array[2520] = 32'hFFFFFFF1;
    // rom_array[2521] = 32'hFFFFFFF0;
    // rom_array[2522] = 32'h00001851;
    // rom_array[2523] = 32'hFFFFFFF0;
    // rom_array[2524] = 32'h00001859;
    // rom_array[2525] = 32'hFFFFFFF0;
    // rom_array[2526] = 32'hFFFFFFF0;
    // rom_array[2527] = 32'hFFFFFFF0;
    // rom_array[2528] = 32'hFFFFFFF0;
    // rom_array[2529] = 32'hFFFFFFF0;
    // rom_array[2530] = 32'h00001861;
    // rom_array[2531] = 32'hFFFFFFF0;
    // rom_array[2532] = 32'h00001869;
    // rom_array[2533] = 32'hFFFFFFF0;
    // rom_array[2534] = 32'h00001871;
    // rom_array[2535] = 32'hFFFFFFF0;
    // rom_array[2536] = 32'hFFFFFFF1;
    // rom_array[2537] = 32'hFFFFFFF0;
    // rom_array[2538] = 32'h00001879;
    // rom_array[2539] = 32'hFFFFFFF0;
    // rom_array[2540] = 32'hFFFFFFF1;
    // rom_array[2541] = 32'hFFFFFFF0;
    // rom_array[2542] = 32'h00001881;
    // rom_array[2543] = 32'hFFFFFFF0;
    // rom_array[2544] = 32'h00001889;
    // rom_array[2545] = 32'hFFFFFFF0;
    // rom_array[2546] = 32'h00001891;
    // rom_array[2547] = 32'hFFFFFFF0;
    // rom_array[2548] = 32'h00001899;
    // rom_array[2549] = 32'hFFFFFFF0;
    // rom_array[2550] = 32'hFFFFFFF0;
    // rom_array[2551] = 32'hFFFFFFF0;
    // rom_array[2552] = 32'h000018a1;
    // rom_array[2553] = 32'hFFFFFFF0;
    // rom_array[2554] = 32'hFFFFFFF0;
    // rom_array[2555] = 32'hFFFFFFF0;
    // rom_array[2556] = 32'hFFFFFFF0;
    // rom_array[2557] = 32'hFFFFFFF0;
    // rom_array[2558] = 32'h000018a9;
    // rom_array[2559] = 32'hFFFFFFF0;
    // rom_array[2560] = 32'h000018b1;
    // rom_array[2561] = 32'hFFFFFFF0;
    // rom_array[2562] = 32'h000018b9;
    // rom_array[2563] = 32'hFFFFFFF0;
    // rom_array[2564] = 32'hFFFFFFF1;
    // rom_array[2565] = 32'hFFFFFFF0;
    // rom_array[2566] = 32'h000018c1;
    // rom_array[2567] = 32'hFFFFFFF0;
    // rom_array[2568] = 32'h000018c9;
    // rom_array[2569] = 32'hFFFFFFF0;
    // rom_array[2570] = 32'hFFFFFFF0;
    // rom_array[2571] = 32'hFFFFFFF0;
    // rom_array[2572] = 32'hFFFFFFF0;
    // rom_array[2573] = 32'hFFFFFFF0;
    // rom_array[2574] = 32'h000018d1;
    // rom_array[2575] = 32'hFFFFFFF0;
    // rom_array[2576] = 32'h000018d9;
    // rom_array[2577] = 32'hFFFFFFF0;
    // rom_array[2578] = 32'hFFFFFFF0;
    // rom_array[2579] = 32'hFFFFFFF0;
    // rom_array[2580] = 32'hFFFFFFF0;
    // rom_array[2581] = 32'hFFFFFFF0;
    // rom_array[2582] = 32'h000018e1;
    // rom_array[2583] = 32'hFFFFFFF0;
    // rom_array[2584] = 32'h000018e9;
    // rom_array[2585] = 32'hFFFFFFF0;
    // rom_array[2586] = 32'hFFFFFFF1;
    // rom_array[2587] = 32'hFFFFFFF0;
    // rom_array[2588] = 32'hFFFFFFF1;
    // rom_array[2589] = 32'hFFFFFFF0;
    // rom_array[2590] = 32'h000018f1;
    // rom_array[2591] = 32'hFFFFFFF0;
    // rom_array[2592] = 32'h000018f9;
    // rom_array[2593] = 32'hFFFFFFF0;
    // rom_array[2594] = 32'hFFFFFFF1;
    // rom_array[2595] = 32'hFFFFFFF0;
    // rom_array[2596] = 32'hFFFFFFF1;
    // rom_array[2597] = 32'hFFFFFFF0;
    // rom_array[2598] = 32'h00001901;
    // rom_array[2599] = 32'hFFFFFFF0;
    // rom_array[2600] = 32'h00001909;
    // rom_array[2601] = 32'hFFFFFFF0;
    // rom_array[2602] = 32'h00001911;
    // rom_array[2603] = 32'hFFFFFFF0;
    // rom_array[2604] = 32'hFFFFFFF1;
    // rom_array[2605] = 32'hFFFFFFF0;
    // rom_array[2606] = 32'h00001919;
    // rom_array[2607] = 32'hFFFFFFF0;
    // rom_array[2608] = 32'hFFFFFFF1;
    // rom_array[2609] = 32'hFFFFFFF0;
    // rom_array[2610] = 32'h00001921;
    // rom_array[2611] = 32'hFFFFFFF0;
    // rom_array[2612] = 32'hFFFFFFF1;
    // rom_array[2613] = 32'hFFFFFFF0;
    // rom_array[2614] = 32'h00001929;
    // rom_array[2615] = 32'hFFFFFFF0;
    // rom_array[2616] = 32'hFFFFFFF1;
    // rom_array[2617] = 32'hFFFFFFF0;
    // rom_array[2618] = 32'h00001931;
    // rom_array[2619] = 32'hFFFFFFF0;
    // rom_array[2620] = 32'hFFFFFFF0;
    // rom_array[2621] = 32'hFFFFFFF0;
    // rom_array[2622] = 32'h00001939;
    // rom_array[2623] = 32'hFFFFFFF0;
    // rom_array[2624] = 32'hFFFFFFF0;
    // rom_array[2625] = 32'hFFFFFFF0;
    // rom_array[2626] = 32'h00001941;
    // rom_array[2627] = 32'hFFFFFFF0;
    // rom_array[2628] = 32'hFFFFFFF1;
    // rom_array[2629] = 32'hFFFFFFF0;
    // rom_array[2630] = 32'h00001949;
    // rom_array[2631] = 32'hFFFFFFF0;
    // rom_array[2632] = 32'hFFFFFFF1;
    // rom_array[2633] = 32'hFFFFFFF0;
    // rom_array[2634] = 32'h00001951;
    // rom_array[2635] = 32'hFFFFFFF0;
    // rom_array[2636] = 32'hFFFFFFF0;
    // rom_array[2637] = 32'hFFFFFFF0;
    // rom_array[2638] = 32'h00001959;
    // rom_array[2639] = 32'hFFFFFFF0;
    // rom_array[2640] = 32'hFFFFFFF0;
    // rom_array[2641] = 32'hFFFFFFF0;
    // rom_array[2642] = 32'h00001961;
    // rom_array[2643] = 32'hFFFFFFF0;
    // rom_array[2644] = 32'hFFFFFFF1;
    // rom_array[2645] = 32'hFFFFFFF0;
    // rom_array[2646] = 32'h00001969;
    // rom_array[2647] = 32'hFFFFFFF0;
    // rom_array[2648] = 32'hFFFFFFF1;
    // rom_array[2649] = 32'h00001971;
    // rom_array[2650] = 32'hFFFFFFF0;
    // rom_array[2651] = 32'h00001979;
    // rom_array[2652] = 32'hFFFFFFF0;
    // rom_array[2653] = 32'h00001981;
    // rom_array[2654] = 32'hFFFFFFF0;
    // rom_array[2655] = 32'hFFFFFFF1;
    // rom_array[2656] = 32'hFFFFFFF0;
    // rom_array[2657] = 32'h00001989;
    // rom_array[2658] = 32'hFFFFFFF0;
    // rom_array[2659] = 32'hFFFFFFF0;
    // rom_array[2660] = 32'hFFFFFFF0;
    // rom_array[2661] = 32'h00001991;
    // rom_array[2662] = 32'hFFFFFFF0;
    // rom_array[2663] = 32'hFFFFFFF0;
    // rom_array[2664] = 32'hFFFFFFF0;
    // rom_array[2665] = 32'h00001999;
    // rom_array[2666] = 32'hFFFFFFF0;
    // rom_array[2667] = 32'hFFFFFFF1;
    // rom_array[2668] = 32'hFFFFFFF0;
    // rom_array[2669] = 32'h000019a1;
    // rom_array[2670] = 32'hFFFFFFF0;
    // rom_array[2671] = 32'hFFFFFFF1;
    // rom_array[2672] = 32'hFFFFFFF0;
    // rom_array[2673] = 32'h000019a9;
    // rom_array[2674] = 32'hFFFFFFF0;
    // rom_array[2675] = 32'hFFFFFFF1;
    // rom_array[2676] = 32'hFFFFFFF0;
    // rom_array[2677] = 32'h000019b1;
    // rom_array[2678] = 32'hFFFFFFF0;
    // rom_array[2679] = 32'hFFFFFFF1;
    // rom_array[2680] = 32'hFFFFFFF0;
    // rom_array[2681] = 32'h000019b9;
    // rom_array[2682] = 32'hFFFFFFF0;
    // rom_array[2683] = 32'hFFFFFFF0;
    // rom_array[2684] = 32'hFFFFFFF0;
    // rom_array[2685] = 32'h000019c1;
    // rom_array[2686] = 32'hFFFFFFF0;
    // rom_array[2687] = 32'h000019c9;
    // rom_array[2688] = 32'hFFFFFFF0;
    // rom_array[2689] = 32'hFFFFFFF0;
    // rom_array[2690] = 32'hFFFFFFF0;
    // rom_array[2691] = 32'hFFFFFFF0;
    // rom_array[2692] = 32'hFFFFFFF0;
    // rom_array[2693] = 32'h000019d1;
    // rom_array[2694] = 32'hFFFFFFF0;
    // rom_array[2695] = 32'h000019d9;
    // rom_array[2696] = 32'hFFFFFFF0;
    // rom_array[2697] = 32'h000019e1;
    // rom_array[2698] = 32'hFFFFFFF0;
    // rom_array[2699] = 32'hFFFFFFF1;
    // rom_array[2700] = 32'hFFFFFFF0;
    // rom_array[2701] = 32'h000019e9;
    // rom_array[2702] = 32'hFFFFFFF0;
    // rom_array[2703] = 32'h000019f1;
    // rom_array[2704] = 32'hFFFFFFF0;
    // rom_array[2705] = 32'hFFFFFFF1;
    // rom_array[2706] = 32'hFFFFFFF0;
    // rom_array[2707] = 32'hFFFFFFF1;
    // rom_array[2708] = 32'hFFFFFFF0;
    // rom_array[2709] = 32'h000019f9;
    // rom_array[2710] = 32'hFFFFFFF0;
    // rom_array[2711] = 32'h00001a01;
    // rom_array[2712] = 32'hFFFFFFF0;
    // rom_array[2713] = 32'h00001a09;
    // rom_array[2714] = 32'hFFFFFFF0;
    // rom_array[2715] = 32'hFFFFFFF1;
    // rom_array[2716] = 32'hFFFFFFF0;
    // rom_array[2717] = 32'h00001a11;
    // rom_array[2718] = 32'hFFFFFFF0;
    // rom_array[2719] = 32'h00001a19;
    // rom_array[2720] = 32'hFFFFFFF0;
    // rom_array[2721] = 32'h00001a21;
    // rom_array[2722] = 32'hFFFFFFF0;
    // rom_array[2723] = 32'hFFFFFFF0;
    // rom_array[2724] = 32'hFFFFFFF0;
    // rom_array[2725] = 32'h00001a29;
    // rom_array[2726] = 32'hFFFFFFF0;
    // rom_array[2727] = 32'hFFFFFFF0;
    // rom_array[2728] = 32'hFFFFFFF0;
    // rom_array[2729] = 32'hFFFFFFF0;
    // rom_array[2730] = 32'hFFFFFFF0;
    // rom_array[2731] = 32'hFFFFFFF0;
    // rom_array[2732] = 32'hFFFFFFF0;
    // rom_array[2733] = 32'h00001a31;
    // rom_array[2734] = 32'hFFFFFFF0;
    // rom_array[2735] = 32'h00001a39;
    // rom_array[2736] = 32'hFFFFFFF0;
    // rom_array[2737] = 32'hFFFFFFF0;
    // rom_array[2738] = 32'hFFFFFFF0;
    // rom_array[2739] = 32'hFFFFFFF0;
    // rom_array[2740] = 32'hFFFFFFF0;
    // rom_array[2741] = 32'h00001a41;
    // rom_array[2742] = 32'hFFFFFFF0;
    // rom_array[2743] = 32'h00001a49;
    // rom_array[2744] = 32'hFFFFFFF0;
    // rom_array[2745] = 32'hFFFFFFF0;
    // rom_array[2746] = 32'hFFFFFFF0;
    // rom_array[2747] = 32'hFFFFFFF0;
    // rom_array[2748] = 32'hFFFFFFF0;
    // rom_array[2749] = 32'h00001a51;
    // rom_array[2750] = 32'hFFFFFFF0;
    // rom_array[2751] = 32'h00001a59;
    // rom_array[2752] = 32'hFFFFFFF0;
    // rom_array[2753] = 32'h00001a61;
    // rom_array[2754] = 32'hFFFFFFF0;
    // rom_array[2755] = 32'hFFFFFFF1;
    // rom_array[2756] = 32'hFFFFFFF0;
    // rom_array[2757] = 32'h00001a69;
    // rom_array[2758] = 32'hFFFFFFF0;
    // rom_array[2759] = 32'h00001a71;
    // rom_array[2760] = 32'hFFFFFFF0;
    // rom_array[2761] = 32'hFFFFFFF1;
    // rom_array[2762] = 32'hFFFFFFF0;
    // rom_array[2763] = 32'h00001a79;
    // rom_array[2764] = 32'hFFFFFFF0;
    // rom_array[2765] = 32'h00001a81;
    // rom_array[2766] = 32'hFFFFFFF0;
    // rom_array[2767] = 32'h00001a89;
    // rom_array[2768] = 32'hFFFFFFF0;
    // rom_array[2769] = 32'hFFFFFFF1;
    // rom_array[2770] = 32'hFFFFFFF0;
    // rom_array[2771] = 32'hFFFFFFF1;
    // rom_array[2772] = 32'hFFFFFFF0;
    // rom_array[2773] = 32'h00001a91;
    // rom_array[2774] = 32'hFFFFFFF0;
    // rom_array[2775] = 32'h00001a99;
    // rom_array[2776] = 32'hFFFFFFF0;
    // rom_array[2777] = 32'hFFFFFFF0;
    // rom_array[2778] = 32'hFFFFFFF0;
    // rom_array[2779] = 32'h00001aa1;
    // rom_array[2780] = 32'hFFFFFFF0;
    // rom_array[2781] = 32'hFFFFFFF0;
    // rom_array[2782] = 32'hFFFFFFF0;
    // rom_array[2783] = 32'h00001aa9;
    // rom_array[2784] = 32'hFFFFFFF0;
    // rom_array[2785] = 32'hFFFFFFF1;
    // rom_array[2786] = 32'hFFFFFFF0;
    // rom_array[2787] = 32'hFFFFFFF1;
    // rom_array[2788] = 32'hFFFFFFF0;
    // rom_array[2789] = 32'h00001ab1;
    // rom_array[2790] = 32'hFFFFFFF0;
    // rom_array[2791] = 32'h00001ab9;
    // rom_array[2792] = 32'hFFFFFFF0;
    // rom_array[2793] = 32'hFFFFFFF0;
    // rom_array[2794] = 32'hFFFFFFF0;
    // rom_array[2795] = 32'h00001ac1;
    // rom_array[2796] = 32'hFFFFFFF0;
    // rom_array[2797] = 32'hFFFFFFF0;
    // rom_array[2798] = 32'hFFFFFFF0;
    // rom_array[2799] = 32'h00001ac9;
    // rom_array[2800] = 32'hFFFFFFF0;
    // rom_array[2801] = 32'h00001ad1;
    // rom_array[2802] = 32'hFFFFFFF0;
    // rom_array[2803] = 32'h00001ad9;
    // rom_array[2804] = 32'hFFFFFFF0;
    // rom_array[2805] = 32'h00001ae1;
    // rom_array[2806] = 32'hFFFFFFF0;
    // rom_array[2807] = 32'h00001ae9;
    // rom_array[2808] = 32'hFFFFFFF0;
    // rom_array[2809] = 32'hFFFFFFF0;
    // rom_array[2810] = 32'hFFFFFFF0;
    // rom_array[2811] = 32'h00001af1;
    // rom_array[2812] = 32'hFFFFFFF0;
    // rom_array[2813] = 32'hFFFFFFF0;
    // rom_array[2814] = 32'hFFFFFFF0;
    // rom_array[2815] = 32'h00001af9;
    // rom_array[2816] = 32'hFFFFFFF0;
    // rom_array[2817] = 32'hFFFFFFF1;
    // rom_array[2818] = 32'hFFFFFFF0;
    // rom_array[2819] = 32'hFFFFFFF1;
    // rom_array[2820] = 32'hFFFFFFF0;
    // rom_array[2821] = 32'hFFFFFFF1;
    // rom_array[2822] = 32'hFFFFFFF0;
    // rom_array[2823] = 32'hFFFFFFF1;
    // rom_array[2824] = 32'hFFFFFFF0;
    // rom_array[2825] = 32'h00001b01;
    // rom_array[2826] = 32'hFFFFFFF0;
    // rom_array[2827] = 32'h00001b09;
    // rom_array[2828] = 32'hFFFFFFF0;
    // rom_array[2829] = 32'h00001b11;
    // rom_array[2830] = 32'hFFFFFFF0;
    // rom_array[2831] = 32'hFFFFFFF1;
    // rom_array[2832] = 32'hFFFFFFF0;
    // rom_array[2833] = 32'h00001b19;
    // rom_array[2834] = 32'hFFFFFFF0;
    // rom_array[2835] = 32'h00001b21;
    // rom_array[2836] = 32'hFFFFFFF0;
    // rom_array[2837] = 32'hFFFFFFF0;
    // rom_array[2838] = 32'hFFFFFFF0;
    // rom_array[2839] = 32'hFFFFFFF0;
    // rom_array[2840] = 32'hFFFFFFF0;
    // rom_array[2841] = 32'h00001b29;
    // rom_array[2842] = 32'hFFFFFFF0;
    // rom_array[2843] = 32'h00001b31;
    // rom_array[2844] = 32'hFFFFFFF0;
    // rom_array[2845] = 32'hFFFFFFF1;
    // rom_array[2846] = 32'hFFFFFFF0;
    // rom_array[2847] = 32'h00001b39;
    // rom_array[2848] = 32'hFFFFFFF0;
    // rom_array[2849] = 32'h00001b41;
    // rom_array[2850] = 32'hFFFFFFF0;
    // rom_array[2851] = 32'h00001b49;
    // rom_array[2852] = 32'hFFFFFFF0;
    // rom_array[2853] = 32'h00001b51;
    // rom_array[2854] = 32'hFFFFFFF0;
    // rom_array[2855] = 32'h00001b59;
    // rom_array[2856] = 32'hFFFFFFF0;
    // rom_array[2857] = 32'h00001b61;
    // rom_array[2858] = 32'hFFFFFFF0;
    // rom_array[2859] = 32'h00001b69;
    // rom_array[2860] = 32'hFFFFFFF0;
    // rom_array[2861] = 32'hFFFFFFF0;
    // rom_array[2862] = 32'hFFFFFFF0;
    // rom_array[2863] = 32'hFFFFFFF0;
    // rom_array[2864] = 32'hFFFFFFF0;
    // rom_array[2865] = 32'h00001b71;
    // rom_array[2866] = 32'hFFFFFFF0;
    // rom_array[2867] = 32'h00001b79;
    // rom_array[2868] = 32'hFFFFFFF0;
    // rom_array[2869] = 32'hFFFFFFF0;
    // rom_array[2870] = 32'hFFFFFFF0;
    // rom_array[2871] = 32'hFFFFFFF0;
    // rom_array[2872] = 32'hFFFFFFF0;
    // rom_array[2873] = 32'h00001b81;
    // rom_array[2874] = 32'hFFFFFFF0;
    // rom_array[2875] = 32'h00001b89;
    // rom_array[2876] = 32'hFFFFFFF0;
    // rom_array[2877] = 32'h00001b91;
    // rom_array[2878] = 32'hFFFFFFF0;
    // rom_array[2879] = 32'hFFFFFFF1;
    // rom_array[2880] = 32'hFFFFFFF0;
    // rom_array[2881] = 32'h00001b99;
    // rom_array[2882] = 32'hFFFFFFF0;
    // rom_array[2883] = 32'h00001ba1;
    // rom_array[2884] = 32'hFFFFFFF0;
    // rom_array[2885] = 32'hFFFFFFF0;
    // rom_array[2886] = 32'hFFFFFFF0;
    // rom_array[2887] = 32'hFFFFFFF0;
    // rom_array[2888] = 32'hFFFFFFF0;
    // rom_array[2889] = 32'h00001ba9;
    // rom_array[2890] = 32'hFFFFFFF0;
    // rom_array[2891] = 32'h00001bb1;
    // rom_array[2892] = 32'hFFFFFFF0;
    // rom_array[2893] = 32'hFFFFFFF1;
    // rom_array[2894] = 32'hFFFFFFF0;
    // rom_array[2895] = 32'hFFFFFFF1;
    // rom_array[2896] = 32'hFFFFFFF0;
    // rom_array[2897] = 32'h00001bb9;
    // rom_array[2898] = 32'hFFFFFFF0;
    // rom_array[2899] = 32'h00001bc1;
    // rom_array[2900] = 32'hFFFFFFF0;
    // rom_array[2901] = 32'hFFFFFFF1;
    // rom_array[2902] = 32'hFFFFFFF0;
    // rom_array[2903] = 32'hFFFFFFF1;
    // rom_array[2904] = 32'hFFFFFFF0;
    // rom_array[2905] = 32'h00001bc9;
    // rom_array[2906] = 32'hFFFFFFF0;
    // rom_array[2907] = 32'h00001bd1;
    // rom_array[2908] = 32'hFFFFFFF0;
    // rom_array[2909] = 32'hFFFFFFF0;
    // rom_array[2910] = 32'hFFFFFFF0;
    // rom_array[2911] = 32'hFFFFFFF0;
    // rom_array[2912] = 32'hFFFFFFF0;
    // rom_array[2913] = 32'h00001bd9;
    // rom_array[2914] = 32'hFFFFFFF0;
    // rom_array[2915] = 32'h00001be1;
    // rom_array[2916] = 32'hFFFFFFF0;
    // rom_array[2917] = 32'h00001be9;
    // rom_array[2918] = 32'hFFFFFFF0;
    // rom_array[2919] = 32'hFFFFFFF1;
    // rom_array[2920] = 32'hFFFFFFF0;
    // rom_array[2921] = 32'h00001bf1;
    // rom_array[2922] = 32'hFFFFFFF0;
    // rom_array[2923] = 32'hFFFFFFF1;
    // rom_array[2924] = 32'hFFFFFFF0;
    // rom_array[2925] = 32'h00001bf9;
    // rom_array[2926] = 32'hFFFFFFF0;
    // rom_array[2927] = 32'h00001c01;
    // rom_array[2928] = 32'hFFFFFFF0;
    // rom_array[2929] = 32'h00001c09;
    // rom_array[2930] = 32'hFFFFFFF0;
    // rom_array[2931] = 32'h00001c11;
    // rom_array[2932] = 32'hFFFFFFF0;
    // rom_array[2933] = 32'hFFFFFFF0;
    // rom_array[2934] = 32'hFFFFFFF0;
    // rom_array[2935] = 32'h00001c19;
    // rom_array[2936] = 32'hFFFFFFF0;
    // rom_array[2937] = 32'hFFFFFFF0;
    // rom_array[2938] = 32'hFFFFFFF0;
    // rom_array[2939] = 32'hFFFFFFF0;
    // rom_array[2940] = 32'hFFFFFFF0;
    // rom_array[2941] = 32'h00001c21;
    // rom_array[2942] = 32'hFFFFFFF0;
    // rom_array[2943] = 32'h00001c29;
    // rom_array[2944] = 32'hFFFFFFF0;
    // rom_array[2945] = 32'h00001c31;
    // rom_array[2946] = 32'hFFFFFFF0;
    // rom_array[2947] = 32'hFFFFFFF1;
    // rom_array[2948] = 32'hFFFFFFF0;
    // rom_array[2949] = 32'h00001c39;
    // rom_array[2950] = 32'hFFFFFFF0;
    // rom_array[2951] = 32'h00001c41;
    // rom_array[2952] = 32'hFFFFFFF0;
    // rom_array[2953] = 32'hFFFFFFF0;
    // rom_array[2954] = 32'hFFFFFFF0;
    // rom_array[2955] = 32'hFFFFFFF0;
    // rom_array[2956] = 32'hFFFFFFF0;
    // rom_array[2957] = 32'h00001c49;
    // rom_array[2958] = 32'hFFFFFFF0;
    // rom_array[2959] = 32'h00001c51;
    // rom_array[2960] = 32'hFFFFFFF0;
    // rom_array[2961] = 32'hFFFFFFF0;
    // rom_array[2962] = 32'hFFFFFFF0;
    // rom_array[2963] = 32'hFFFFFFF0;
    // rom_array[2964] = 32'hFFFFFFF0;
    // rom_array[2965] = 32'h00001c59;
    // rom_array[2966] = 32'hFFFFFFF0;
    // rom_array[2967] = 32'h00001c61;
    // rom_array[2968] = 32'hFFFFFFF0;
    // rom_array[2969] = 32'hFFFFFFF1;
    // rom_array[2970] = 32'hFFFFFFF0;
    // rom_array[2971] = 32'hFFFFFFF1;
    // rom_array[2972] = 32'hFFFFFFF0;
    // rom_array[2973] = 32'h00001c69;
    // rom_array[2974] = 32'hFFFFFFF0;
    // rom_array[2975] = 32'h00001c71;
    // rom_array[2976] = 32'hFFFFFFF0;
    // rom_array[2977] = 32'hFFFFFFF1;
    // rom_array[2978] = 32'hFFFFFFF0;
    // rom_array[2979] = 32'hFFFFFFF1;
    // rom_array[2980] = 32'hFFFFFFF0;
    // rom_array[2981] = 32'h00001c79;
    // rom_array[2982] = 32'hFFFFFFF0;
    // rom_array[2983] = 32'h00001c81;
    // rom_array[2984] = 32'hFFFFFFF0;
    // rom_array[2985] = 32'h00001c89;
    // rom_array[2986] = 32'hFFFFFFF0;
    // rom_array[2987] = 32'hFFFFFFF1;
    // rom_array[2988] = 32'hFFFFFFF0;
    // rom_array[2989] = 32'h00001c91;
    // rom_array[2990] = 32'hFFFFFFF0;
    // rom_array[2991] = 32'hFFFFFFF1;
    // rom_array[2992] = 32'hFFFFFFF0;
    // rom_array[2993] = 32'h00001c99;
    // rom_array[2994] = 32'hFFFFFFF0;
    // rom_array[2995] = 32'hFFFFFFF1;
    // rom_array[2996] = 32'hFFFFFFF0;
    // rom_array[2997] = 32'h00001ca1;
    // rom_array[2998] = 32'hFFFFFFF0;
    // rom_array[2999] = 32'hFFFFFFF1;
    // rom_array[3000] = 32'hFFFFFFF0;
    // rom_array[3001] = 32'h00001ca9;
    // rom_array[3002] = 32'hFFFFFFF0;
    // rom_array[3003] = 32'hFFFFFFF0;
    // rom_array[3004] = 32'hFFFFFFF0;
    // rom_array[3005] = 32'h00001cb1;
    // rom_array[3006] = 32'hFFFFFFF0;
    // rom_array[3007] = 32'hFFFFFFF0;
    // rom_array[3008] = 32'hFFFFFFF0;
    // rom_array[3009] = 32'h00001cb9;
    // rom_array[3010] = 32'hFFFFFFF0;
    // rom_array[3011] = 32'hFFFFFFF1;
    // rom_array[3012] = 32'hFFFFFFF0;
    // rom_array[3013] = 32'h00001cc1;
    // rom_array[3014] = 32'hFFFFFFF0;
    // rom_array[3015] = 32'hFFFFFFF1;
    // rom_array[3016] = 32'hFFFFFFF0;
    // rom_array[3017] = 32'h00001cc9;
    // rom_array[3018] = 32'hFFFFFFF0;
    // rom_array[3019] = 32'hFFFFFFF0;
    // rom_array[3020] = 32'hFFFFFFF0;
    // rom_array[3021] = 32'h00001cd1;
    // rom_array[3022] = 32'hFFFFFFF0;
    // rom_array[3023] = 32'hFFFFFFF0;
    // rom_array[3024] = 32'hFFFFFFF0;
    // rom_array[3025] = 32'h00001cd9;
    // rom_array[3026] = 32'hFFFFFFF0;
    // rom_array[3027] = 32'hFFFFFFF1;
    // rom_array[3028] = 32'hFFFFFFF0;
    // rom_array[3029] = 32'h00001ce1;
    // rom_array[3030] = 32'hFFFFFFF0;
    // rom_array[3031] = 32'hFFFFFFF1;
    // rom_array[3032] = 32'hFFFFFFF0;
    // rom_array[3033] = 32'hFFFFFFF0;
    // rom_array[3034] = 32'hFFFFFFF0;
    // rom_array[3035] = 32'hFFFFFFF0;
    // rom_array[3036] = 32'h00001ce9;
    // rom_array[3037] = 32'hFFFFFFF0;
    // rom_array[3038] = 32'hFFFFFFF0;
    // rom_array[3039] = 32'hFFFFFFF0;
    // rom_array[3040] = 32'h00001cf1;
    // rom_array[3041] = 32'hFFFFFFF0;
    // rom_array[3042] = 32'h00001cf9;
    // rom_array[3043] = 32'hFFFFFFF0;
    // rom_array[3044] = 32'h00001d01;
    // rom_array[3045] = 32'hFFFFFFF0;
    // rom_array[3046] = 32'hFFFFFFF1;
    // rom_array[3047] = 32'hFFFFFFF0;
    // rom_array[3048] = 32'h00001d09;
    // rom_array[3049] = 32'hFFFFFFF0;
    // rom_array[3050] = 32'hFFFFFFF0;
    // rom_array[3051] = 32'hFFFFFFF0;
    // rom_array[3052] = 32'hFFFFFFF0;
    // rom_array[3053] = 32'hFFFFFFF0;
    // rom_array[3054] = 32'h00001d11;
    // rom_array[3055] = 32'hFFFFFFF0;
    // rom_array[3056] = 32'h00001d19;
    // rom_array[3057] = 32'hFFFFFFF0;
    // rom_array[3058] = 32'hFFFFFFF0;
    // rom_array[3059] = 32'hFFFFFFF0;
    // rom_array[3060] = 32'h00001d21;
    // rom_array[3061] = 32'hFFFFFFF0;
    // rom_array[3062] = 32'h00001d29;
    // rom_array[3063] = 32'hFFFFFFF0;
    // rom_array[3064] = 32'h00001d31;
    // rom_array[3065] = 32'hFFFFFFF0;
    // rom_array[3066] = 32'hFFFFFFF1;
    // rom_array[3067] = 32'hFFFFFFF0;
    // rom_array[3068] = 32'hFFFFFFF1;
    // rom_array[3069] = 32'hFFFFFFF0;
    // rom_array[3070] = 32'h00001d39;
    // rom_array[3071] = 32'hFFFFFFF0;
    // rom_array[3072] = 32'h00001d41;
    // rom_array[3073] = 32'hFFFFFFF0;
    // rom_array[3074] = 32'hFFFFFFF1;
    // rom_array[3075] = 32'hFFFFFFF0;
    // rom_array[3076] = 32'h00001d49;
    // rom_array[3077] = 32'hFFFFFFF0;
    // rom_array[3078] = 32'h00001d51;
    // rom_array[3079] = 32'hFFFFFFF0;
    // rom_array[3080] = 32'h00001d59;
    // rom_array[3081] = 32'hFFFFFFF0;
    // rom_array[3082] = 32'hFFFFFFF1;
    // rom_array[3083] = 32'hFFFFFFF0;
    // rom_array[3084] = 32'h00001d61;
    // rom_array[3085] = 32'hFFFFFFF0;
    // rom_array[3086] = 32'hFFFFFFF1;
    // rom_array[3087] = 32'hFFFFFFF0;
    // rom_array[3088] = 32'h00001d69;
    // rom_array[3089] = 32'hFFFFFFF0;
    // rom_array[3090] = 32'hFFFFFFF1;
    // rom_array[3091] = 32'hFFFFFFF0;
    // rom_array[3092] = 32'h00001d71;
    // rom_array[3093] = 32'hFFFFFFF0;
    // rom_array[3094] = 32'hFFFFFFF1;
    // rom_array[3095] = 32'hFFFFFFF0;
    // rom_array[3096] = 32'h00001d79;
    // rom_array[3097] = 32'hFFFFFFF0;
    // rom_array[3098] = 32'hFFFFFFF0;
    // rom_array[3099] = 32'hFFFFFFF0;
    // rom_array[3100] = 32'h00001d81;
    // rom_array[3101] = 32'hFFFFFFF0;
    // rom_array[3102] = 32'hFFFFFFF0;
    // rom_array[3103] = 32'hFFFFFFF0;
    // rom_array[3104] = 32'h00001d89;
    // rom_array[3105] = 32'hFFFFFFF0;
    // rom_array[3106] = 32'hFFFFFFF1;
    // rom_array[3107] = 32'hFFFFFFF0;
    // rom_array[3108] = 32'h00001d91;
    // rom_array[3109] = 32'hFFFFFFF0;
    // rom_array[3110] = 32'h00001d99;
    // rom_array[3111] = 32'hFFFFFFF0;
    // rom_array[3112] = 32'h00001da1;
    // rom_array[3113] = 32'hFFFFFFF0;
    // rom_array[3114] = 32'hFFFFFFF0;
    // rom_array[3115] = 32'hFFFFFFF0;
    // rom_array[3116] = 32'hFFFFFFF0;
    // rom_array[3117] = 32'hFFFFFFF0;
    // rom_array[3118] = 32'h00001da9;
    // rom_array[3119] = 32'hFFFFFFF0;
    // rom_array[3120] = 32'h00001db1;
    // rom_array[3121] = 32'hFFFFFFF0;
    // rom_array[3122] = 32'hFFFFFFF0;
    // rom_array[3123] = 32'hFFFFFFF0;
    // rom_array[3124] = 32'hFFFFFFF0;
    // rom_array[3125] = 32'hFFFFFFF0;
    // rom_array[3126] = 32'h00001db9;
    // rom_array[3127] = 32'hFFFFFFF0;
    // rom_array[3128] = 32'h00001dc1;
    // rom_array[3129] = 32'hFFFFFFF0;
    // rom_array[3130] = 32'hFFFFFFF0;
    // rom_array[3131] = 32'hFFFFFFF0;
    // rom_array[3132] = 32'hFFFFFFF0;
    // rom_array[3133] = 32'hFFFFFFF0;
    // rom_array[3134] = 32'h00001dc9;
    // rom_array[3135] = 32'hFFFFFFF0;
    // rom_array[3136] = 32'h00001dd1;
    // rom_array[3137] = 32'hFFFFFFF0;
    // rom_array[3138] = 32'hFFFFFFF1;
    // rom_array[3139] = 32'hFFFFFFF0;
    // rom_array[3140] = 32'hFFFFFFF1;
    // rom_array[3141] = 32'hFFFFFFF0;
    // rom_array[3142] = 32'h00001dd9;
    // rom_array[3143] = 32'hFFFFFFF0;
    // rom_array[3144] = 32'h00001de1;
    // rom_array[3145] = 32'hFFFFFFF0;
    // rom_array[3146] = 32'hFFFFFFF1;
    // rom_array[3147] = 32'hFFFFFFF0;
    // rom_array[3148] = 32'hFFFFFFF1;
    // rom_array[3149] = 32'hFFFFFFF0;
    // rom_array[3150] = 32'h00001de9;
    // rom_array[3151] = 32'hFFFFFFF0;
    // rom_array[3152] = 32'h00001df1;
    // rom_array[3153] = 32'hFFFFFFF0;
    // rom_array[3154] = 32'hFFFFFFF1;
    // rom_array[3155] = 32'hFFFFFFF0;
    // rom_array[3156] = 32'hFFFFFFF1;
    // rom_array[3157] = 32'hFFFFFFF0;
    // rom_array[3158] = 32'hFFFFFFF1;
    // rom_array[3159] = 32'hFFFFFFF0;
    // rom_array[3160] = 32'hFFFFFFF1;
    // rom_array[3161] = 32'hFFFFFFF0;
    // rom_array[3162] = 32'hFFFFFFF1;
    // rom_array[3163] = 32'hFFFFFFF0;
    // rom_array[3164] = 32'hFFFFFFF1;
    // rom_array[3165] = 32'hFFFFFFF0;
    // rom_array[3166] = 32'hFFFFFFF1;
    // rom_array[3167] = 32'hFFFFFFF0;
    // rom_array[3168] = 32'hFFFFFFF1;
    // rom_array[3169] = 32'hFFFFFFF0;
    // rom_array[3170] = 32'hFFFFFFF1;
    // rom_array[3171] = 32'hFFFFFFF0;
    // rom_array[3172] = 32'h00001df9;
    // rom_array[3173] = 32'hFFFFFFF0;
    // rom_array[3174] = 32'h00001e01;
    // rom_array[3175] = 32'hFFFFFFF0;
    // rom_array[3176] = 32'h00001e09;
    // rom_array[3177] = 32'hFFFFFFF0;
    // rom_array[3178] = 32'hFFFFFFF1;
    // rom_array[3179] = 32'hFFFFFFF0;
    // rom_array[3180] = 32'h00001e11;
    // rom_array[3181] = 32'hFFFFFFF0;
    // rom_array[3182] = 32'hFFFFFFF1;
    // rom_array[3183] = 32'hFFFFFFF0;
    // rom_array[3184] = 32'h00001e19;
    // rom_array[3185] = 32'hFFFFFFF0;
    // rom_array[3186] = 32'h00001e21;
    // rom_array[3187] = 32'hFFFFFFF0;
    // rom_array[3188] = 32'h00001e29;
    // rom_array[3189] = 32'hFFFFFFF0;
    // rom_array[3190] = 32'h00001e31;
    // rom_array[3191] = 32'hFFFFFFF0;
    // rom_array[3192] = 32'h00001e39;
    // rom_array[3193] = 32'hFFFFFFF0;
    // rom_array[3194] = 32'h00001e41;
    // rom_array[3195] = 32'hFFFFFFF0;
    // rom_array[3196] = 32'h00001e49;
    // rom_array[3197] = 32'hFFFFFFF0;
    // rom_array[3198] = 32'h00001e51;
    // rom_array[3199] = 32'hFFFFFFF0;
    // rom_array[3200] = 32'h00001e59;
    // rom_array[3201] = 32'hFFFFFFF0;
    // rom_array[3202] = 32'hFFFFFFF1;
    // rom_array[3203] = 32'hFFFFFFF0;
    // rom_array[3204] = 32'hFFFFFFF1;
    // rom_array[3205] = 32'hFFFFFFF0;
    // rom_array[3206] = 32'hFFFFFFF1;
    // rom_array[3207] = 32'hFFFFFFF0;
    // rom_array[3208] = 32'hFFFFFFF1;
    // rom_array[3209] = 32'hFFFFFFF0;
    // rom_array[3210] = 32'hFFFFFFF1;
    // rom_array[3211] = 32'hFFFFFFF0;
    // rom_array[3212] = 32'hFFFFFFF1;
    // rom_array[3213] = 32'hFFFFFFF0;
    // rom_array[3214] = 32'hFFFFFFF1;
    // rom_array[3215] = 32'hFFFFFFF0;
    // rom_array[3216] = 32'hFFFFFFF1;
    // rom_array[3217] = 32'hFFFFFFF0;
    // rom_array[3218] = 32'h00001e61;
    // rom_array[3219] = 32'hFFFFFFF0;
    // rom_array[3220] = 32'h00001e69;
    // rom_array[3221] = 32'hFFFFFFF0;
    // rom_array[3222] = 32'h00001e71;
    // rom_array[3223] = 32'hFFFFFFF0;
    // rom_array[3224] = 32'h00001e79;
    // rom_array[3225] = 32'hFFFFFFF0;
    // rom_array[3226] = 32'hFFFFFFF1;
    // rom_array[3227] = 32'hFFFFFFF0;
    // rom_array[3228] = 32'h00001e81;
    // rom_array[3229] = 32'hFFFFFFF0;
    // rom_array[3230] = 32'hFFFFFFF1;
    // rom_array[3231] = 32'hFFFFFFF0;
    // rom_array[3232] = 32'h00001e89;
    // rom_array[3233] = 32'hFFFFFFF0;
    // rom_array[3234] = 32'h00001e91;
    // rom_array[3235] = 32'hFFFFFFF0;
    // rom_array[3236] = 32'h00001e99;
    // rom_array[3237] = 32'hFFFFFFF0;
    // rom_array[3238] = 32'h00001ea1;
    // rom_array[3239] = 32'hFFFFFFF0;
    // rom_array[3240] = 32'h00001ea9;
    // rom_array[3241] = 32'hFFFFFFF0;
    // rom_array[3242] = 32'h00001eb1;
    // rom_array[3243] = 32'hFFFFFFF0;
    // rom_array[3244] = 32'h00001eb9;
    // rom_array[3245] = 32'hFFFFFFF0;
    // rom_array[3246] = 32'h00001ec1;
    // rom_array[3247] = 32'hFFFFFFF0;
    // rom_array[3248] = 32'h00001ec9;
    // rom_array[3249] = 32'hFFFFFFF0;
    // rom_array[3250] = 32'h00001ed1;
    // rom_array[3251] = 32'hFFFFFFF0;
    // rom_array[3252] = 32'h00001ed9;
    // rom_array[3253] = 32'hFFFFFFF0;
    // rom_array[3254] = 32'hFFFFFFF0;
    // rom_array[3255] = 32'hFFFFFFF0;
    // rom_array[3256] = 32'hFFFFFFF0;
    // rom_array[3257] = 32'hFFFFFFF0;
    // rom_array[3258] = 32'h00001ee1;
    // rom_array[3259] = 32'hFFFFFFF0;
    // rom_array[3260] = 32'h00001ee9;
    // rom_array[3261] = 32'hFFFFFFF0;
    // rom_array[3262] = 32'hFFFFFFF0;
    // rom_array[3263] = 32'hFFFFFFF0;
    // rom_array[3264] = 32'hFFFFFFF0;
    // rom_array[3265] = 32'hFFFFFFF0;
    // rom_array[3266] = 32'h00001ef1;
    // rom_array[3267] = 32'hFFFFFFF0;
    // rom_array[3268] = 32'h00001ef9;
    // rom_array[3269] = 32'hFFFFFFF0;
    // rom_array[3270] = 32'h00001f01;
    // rom_array[3271] = 32'hFFFFFFF0;
    // rom_array[3272] = 32'h00001f09;
    // rom_array[3273] = 32'hFFFFFFF0;
    // rom_array[3274] = 32'h00001f11;
    // rom_array[3275] = 32'hFFFFFFF0;
    // rom_array[3276] = 32'h00001f19;
    // rom_array[3277] = 32'hFFFFFFF0;
    // rom_array[3278] = 32'hFFFFFFF0;
    // rom_array[3279] = 32'hFFFFFFF0;
    // rom_array[3280] = 32'hFFFFFFF0;
    // rom_array[3281] = 32'hFFFFFFF0;
    // rom_array[3282] = 32'h00001f21;
    // rom_array[3283] = 32'hFFFFFFF0;
    // rom_array[3284] = 32'h00001f29;
    // rom_array[3285] = 32'hFFFFFFF0;
    // rom_array[3286] = 32'hFFFFFFF1;
    // rom_array[3287] = 32'hFFFFFFF0;
    // rom_array[3288] = 32'hFFFFFFF1;
    // rom_array[3289] = 32'hFFFFFFF0;
    // rom_array[3290] = 32'h00001f31;
    // rom_array[3291] = 32'hFFFFFFF0;
    // rom_array[3292] = 32'h00001f39;
    // rom_array[3293] = 32'hFFFFFFF0;
    // rom_array[3294] = 32'hFFFFFFF1;
    // rom_array[3295] = 32'hFFFFFFF0;
    // rom_array[3296] = 32'hFFFFFFF1;
    // rom_array[3297] = 32'hFFFFFFF0;
    // rom_array[3298] = 32'h00001f41;
    // rom_array[3299] = 32'hFFFFFFF0;
    // rom_array[3300] = 32'h00001f49;
    // rom_array[3301] = 32'hFFFFFFF0;
    // rom_array[3302] = 32'h00001f51;
    // rom_array[3303] = 32'hFFFFFFF0;
    // rom_array[3304] = 32'hFFFFFFF0;
    // rom_array[3305] = 32'hFFFFFFF0;
    // rom_array[3306] = 32'h00001f59;
    // rom_array[3307] = 32'hFFFFFFF0;
    // rom_array[3308] = 32'h00001f61;
    // rom_array[3309] = 32'hFFFFFFF0;
    // rom_array[3310] = 32'hFFFFFFF0;
    // rom_array[3311] = 32'hFFFFFFF0;
    // rom_array[3312] = 32'h00001f69;
    // rom_array[3313] = 32'hFFFFFFF0;
    // rom_array[3314] = 32'h00001f71;
    // rom_array[3315] = 32'hFFFFFFF0;
    // rom_array[3316] = 32'h00001f79;
    // rom_array[3317] = 32'hFFFFFFF0;
    // rom_array[3318] = 32'hFFFFFFF1;
    // rom_array[3319] = 32'hFFFFFFF0;
    // rom_array[3320] = 32'h00001f81;
    // rom_array[3321] = 32'hFFFFFFF0;
    // rom_array[3322] = 32'h00001f89;
    // rom_array[3323] = 32'hFFFFFFF0;
    // rom_array[3324] = 32'h00001f91;
    // rom_array[3325] = 32'hFFFFFFF0;
    // rom_array[3326] = 32'hFFFFFFF1;
    // rom_array[3327] = 32'hFFFFFFF0;
    // rom_array[3328] = 32'h00001f99;
    // rom_array[3329] = 32'hFFFFFFF0;
    // rom_array[3330] = 32'h00001fa1;
    // rom_array[3331] = 32'hFFFFFFF0;
    // rom_array[3332] = 32'hFFFFFFF0;
    // rom_array[3333] = 32'hFFFFFFF0;
    // rom_array[3334] = 32'h00001fa9;
    // rom_array[3335] = 32'hFFFFFFF0;
    // rom_array[3336] = 32'h00001fb1;
    // rom_array[3337] = 32'hFFFFFFF0;
    // rom_array[3338] = 32'hFFFFFFF0;
    // rom_array[3339] = 32'hFFFFFFF0;
    // rom_array[3340] = 32'h00001fb9;
    // rom_array[3341] = 32'hFFFFFFF0;
    // rom_array[3342] = 32'h00001fc1;
    // rom_array[3343] = 32'hFFFFFFF0;
    // rom_array[3344] = 32'h00001fc9;
    // rom_array[3345] = 32'hFFFFFFF0;
    // rom_array[3346] = 32'h00001fd1;
    // rom_array[3347] = 32'hFFFFFFF0;
    // rom_array[3348] = 32'hFFFFFFF1;
    // rom_array[3349] = 32'hFFFFFFF0;
    // rom_array[3350] = 32'h00001fd9;
    // rom_array[3351] = 32'hFFFFFFF0;
    // rom_array[3352] = 32'h00001fe1;
    // rom_array[3353] = 32'hFFFFFFF0;
    // rom_array[3354] = 32'hFFFFFFF1;
    // rom_array[3355] = 32'hFFFFFFF0;
    // rom_array[3356] = 32'h00001fe9;
    // rom_array[3357] = 32'hFFFFFFF0;
    // rom_array[3358] = 32'h00001ff1;
    // rom_array[3359] = 32'hFFFFFFF0;
    // rom_array[3360] = 32'h00001ff9;
    // rom_array[3361] = 32'hFFFFFFF0;
    // rom_array[3362] = 32'hFFFFFFF1;
    // rom_array[3363] = 32'hFFFFFFF0;
    // rom_array[3364] = 32'h00002001;
    // rom_array[3365] = 32'hFFFFFFF0;
    // rom_array[3366] = 32'hFFFFFFF1;
    // rom_array[3367] = 32'hFFFFFFF0;
    // rom_array[3368] = 32'h00002009;
    // rom_array[3369] = 32'hFFFFFFF0;
    // rom_array[3370] = 32'h00002011;
    // rom_array[3371] = 32'hFFFFFFF0;
    // rom_array[3372] = 32'h00002019;
    // rom_array[3373] = 32'hFFFFFFF0;
    // rom_array[3374] = 32'hFFFFFFF0;
    // rom_array[3375] = 32'hFFFFFFF0;
    // rom_array[3376] = 32'hFFFFFFF0;
    // rom_array[3377] = 32'hFFFFFFF0;
    // rom_array[3378] = 32'hFFFFFFF0;
    // rom_array[3379] = 32'hFFFFFFF0;
    // rom_array[3380] = 32'hFFFFFFF0;
    // rom_array[3381] = 32'hFFFFFFF0;
    // rom_array[3382] = 32'h00002021;
    // rom_array[3383] = 32'hFFFFFFF0;
    // rom_array[3384] = 32'h00002029;
    // rom_array[3385] = 32'hFFFFFFF0;
    // rom_array[3386] = 32'hFFFFFFF0;
    // rom_array[3387] = 32'hFFFFFFF0;
    // rom_array[3388] = 32'hFFFFFFF0;
    // rom_array[3389] = 32'hFFFFFFF0;
    // rom_array[3390] = 32'h00002031;
    // rom_array[3391] = 32'hFFFFFFF0;
    // rom_array[3392] = 32'h00002039;
    // rom_array[3393] = 32'hFFFFFFF0;
    // rom_array[3394] = 32'hFFFFFFF1;
    // rom_array[3395] = 32'hFFFFFFF0;
    // rom_array[3396] = 32'hFFFFFFF1;
    // rom_array[3397] = 32'hFFFFFFF0;
    // rom_array[3398] = 32'h00002041;
    // rom_array[3399] = 32'hFFFFFFF0;
    // rom_array[3400] = 32'h00002049;
    // rom_array[3401] = 32'hFFFFFFF0;
    // rom_array[3402] = 32'hFFFFFFF1;
    // rom_array[3403] = 32'hFFFFFFF0;
    // rom_array[3404] = 32'hFFFFFFF1;
    // rom_array[3405] = 32'hFFFFFFF0;
    // rom_array[3406] = 32'h00002051;
    // rom_array[3407] = 32'hFFFFFFF0;
    // rom_array[3408] = 32'h00002059;
    // rom_array[3409] = 32'hFFFFFFF0;
    // rom_array[3410] = 32'hFFFFFFF0;
    // rom_array[3411] = 32'hFFFFFFF0;
    // rom_array[3412] = 32'hFFFFFFF0;
    // rom_array[3413] = 32'hFFFFFFF0;
    // rom_array[3414] = 32'h00002061;
    // rom_array[3415] = 32'hFFFFFFF0;
    // rom_array[3416] = 32'h00002069;
    // rom_array[3417] = 32'hFFFFFFF0;
    // rom_array[3418] = 32'hFFFFFFF1;
    // rom_array[3419] = 32'hFFFFFFF0;
    // rom_array[3420] = 32'h00002071;
    // rom_array[3421] = 32'hFFFFFFF0;
    // rom_array[3422] = 32'h00002079;
    // rom_array[3423] = 32'hFFFFFFF0;
    // rom_array[3424] = 32'h00002081;
    // rom_array[3425] = 32'hFFFFFFF0;
    // rom_array[3426] = 32'h00002089;
    // rom_array[3427] = 32'hFFFFFFF0;
    // rom_array[3428] = 32'hFFFFFFF0;
    // rom_array[3429] = 32'hFFFFFFF0;
    // rom_array[3430] = 32'h00002091;
    // rom_array[3431] = 32'hFFFFFFF0;
    // rom_array[3432] = 32'hFFFFFFF0;
    // rom_array[3433] = 32'hFFFFFFF0;
    // rom_array[3434] = 32'hFFFFFFF0;
    // rom_array[3435] = 32'hFFFFFFF0;
    // rom_array[3436] = 32'h00002099;
    // rom_array[3437] = 32'hFFFFFFF0;
    // rom_array[3438] = 32'hFFFFFFF0;
    // rom_array[3439] = 32'hFFFFFFF0;
    // rom_array[3440] = 32'h000020a1;
    // rom_array[3441] = 32'hFFFFFFF0;
    // rom_array[3442] = 32'h000020a9;
    // rom_array[3443] = 32'hFFFFFFF0;
    // rom_array[3444] = 32'hFFFFFFF0;
    // rom_array[3445] = 32'hFFFFFFF0;
    // rom_array[3446] = 32'h000020b1;
    // rom_array[3447] = 32'hFFFFFFF0;
    // rom_array[3448] = 32'hFFFFFFF0;
    // rom_array[3449] = 32'hFFFFFFF0;
    // rom_array[3450] = 32'hFFFFFFF0;
    // rom_array[3451] = 32'hFFFFFFF0;
    // rom_array[3452] = 32'h000020b9;
    // rom_array[3453] = 32'hFFFFFFF0;
    // rom_array[3454] = 32'hFFFFFFF0;
    // rom_array[3455] = 32'hFFFFFFF0;
    // rom_array[3456] = 32'h000020c1;
    // rom_array[3457] = 32'hFFFFFFF0;
    // rom_array[3458] = 32'hFFFFFFF1;
    // rom_array[3459] = 32'hFFFFFFF0;
    // rom_array[3460] = 32'h000020c9;
    // rom_array[3461] = 32'hFFFFFFF0;
    // rom_array[3462] = 32'hFFFFFFF1;
    // rom_array[3463] = 32'hFFFFFFF0;
    // rom_array[3464] = 32'h000020d1;
    // rom_array[3465] = 32'hFFFFFFF0;
    // rom_array[3466] = 32'hFFFFFFF1;
    // rom_array[3467] = 32'hFFFFFFF0;
    // rom_array[3468] = 32'h000020d9;
    // rom_array[3469] = 32'hFFFFFFF0;
    // rom_array[3470] = 32'hFFFFFFF1;
    // rom_array[3471] = 32'hFFFFFFF0;
    // rom_array[3472] = 32'h000020e1;
    // rom_array[3473] = 32'hFFFFFFF0;
    // rom_array[3474] = 32'hFFFFFFF0;
    // rom_array[3475] = 32'h000020e9;
    // rom_array[3476] = 32'hFFFFFFF0;
    // rom_array[3477] = 32'hFFFFFFF0;
    // rom_array[3478] = 32'hFFFFFFF0;
    // rom_array[3479] = 32'h000020f1;
    // rom_array[3480] = 32'hFFFFFFF0;
    // rom_array[3481] = 32'h000020f9;
    // rom_array[3482] = 32'hFFFFFFF0;
    // rom_array[3483] = 32'h00002101;
    // rom_array[3484] = 32'hFFFFFFF0;
    // rom_array[3485] = 32'hFFFFFFF1;
    // rom_array[3486] = 32'hFFFFFFF0;
    // rom_array[3487] = 32'h00002109;
    // rom_array[3488] = 32'hFFFFFFF0;
    // rom_array[3489] = 32'hFFFFFFF0;
    // rom_array[3490] = 32'hFFFFFFF0;
    // rom_array[3491] = 32'hFFFFFFF0;
    // rom_array[3492] = 32'hFFFFFFF0;
    // rom_array[3493] = 32'h00002111;
    // rom_array[3494] = 32'hFFFFFFF0;
    // rom_array[3495] = 32'h00002119;
    // rom_array[3496] = 32'hFFFFFFF0;
    // rom_array[3497] = 32'hFFFFFFF0;
    // rom_array[3498] = 32'hFFFFFFF0;
    // rom_array[3499] = 32'h00002121;
    // rom_array[3500] = 32'hFFFFFFF0;
    // rom_array[3501] = 32'h00002129;
    // rom_array[3502] = 32'hFFFFFFF0;
    // rom_array[3503] = 32'h00002131;
    // rom_array[3504] = 32'hFFFFFFF0;
    // rom_array[3505] = 32'hFFFFFFF1;
    // rom_array[3506] = 32'hFFFFFFF0;
    // rom_array[3507] = 32'hFFFFFFF1;
    // rom_array[3508] = 32'hFFFFFFF0;
    // rom_array[3509] = 32'h00002139;
    // rom_array[3510] = 32'hFFFFFFF0;
    // rom_array[3511] = 32'h00002141;
    // rom_array[3512] = 32'hFFFFFFF0;
    // rom_array[3513] = 32'hFFFFFFF1;
    // rom_array[3514] = 32'hFFFFFFF0;
    // rom_array[3515] = 32'h00002149;
    // rom_array[3516] = 32'hFFFFFFF0;
    // rom_array[3517] = 32'h00002151;
    // rom_array[3518] = 32'hFFFFFFF0;
    // rom_array[3519] = 32'h00002159;
    // rom_array[3520] = 32'hFFFFFFF0;
    // rom_array[3521] = 32'hFFFFFFF1;
    // rom_array[3522] = 32'hFFFFFFF0;
    // rom_array[3523] = 32'h00002161;
    // rom_array[3524] = 32'hFFFFFFF0;
    // rom_array[3525] = 32'hFFFFFFF1;
    // rom_array[3526] = 32'hFFFFFFF0;
    // rom_array[3527] = 32'h00002169;
    // rom_array[3528] = 32'hFFFFFFF0;
    // rom_array[3529] = 32'hFFFFFFF1;
    // rom_array[3530] = 32'hFFFFFFF0;
    // rom_array[3531] = 32'h00002171;
    // rom_array[3532] = 32'hFFFFFFF0;
    // rom_array[3533] = 32'hFFFFFFF1;
    // rom_array[3534] = 32'hFFFFFFF0;
    // rom_array[3535] = 32'h00002179;
    // rom_array[3536] = 32'hFFFFFFF0;
    // rom_array[3537] = 32'hFFFFFFF0;
    // rom_array[3538] = 32'hFFFFFFF0;
    // rom_array[3539] = 32'h00002181;
    // rom_array[3540] = 32'hFFFFFFF0;
    // rom_array[3541] = 32'hFFFFFFF0;
    // rom_array[3542] = 32'hFFFFFFF0;
    // rom_array[3543] = 32'h00002189;
    // rom_array[3544] = 32'hFFFFFFF0;
    // rom_array[3545] = 32'hFFFFFFF1;
    // rom_array[3546] = 32'hFFFFFFF0;
    // rom_array[3547] = 32'h00002191;
    // rom_array[3548] = 32'hFFFFFFF0;
    // rom_array[3549] = 32'h00002199;
    // rom_array[3550] = 32'hFFFFFFF0;
    // rom_array[3551] = 32'h000021a1;
    // rom_array[3552] = 32'hFFFFFFF0;
    // rom_array[3553] = 32'hFFFFFFF0;
    // rom_array[3554] = 32'hFFFFFFF0;
    // rom_array[3555] = 32'hFFFFFFF0;
    // rom_array[3556] = 32'hFFFFFFF0;
    // rom_array[3557] = 32'h000021a9;
    // rom_array[3558] = 32'hFFFFFFF0;
    // rom_array[3559] = 32'h000021b1;
    // rom_array[3560] = 32'hFFFFFFF0;
    // rom_array[3561] = 32'hFFFFFFF0;
    // rom_array[3562] = 32'hFFFFFFF0;
    // rom_array[3563] = 32'hFFFFFFF0;
    // rom_array[3564] = 32'hFFFFFFF0;
    // rom_array[3565] = 32'h000021b9;
    // rom_array[3566] = 32'hFFFFFFF0;
    // rom_array[3567] = 32'h000021c1;
    // rom_array[3568] = 32'hFFFFFFF0;
    // rom_array[3569] = 32'hFFFFFFF0;
    // rom_array[3570] = 32'hFFFFFFF0;
    // rom_array[3571] = 32'hFFFFFFF0;
    // rom_array[3572] = 32'hFFFFFFF0;
    // rom_array[3573] = 32'h000021c9;
    // rom_array[3574] = 32'hFFFFFFF0;
    // rom_array[3575] = 32'h000021d1;
    // rom_array[3576] = 32'hFFFFFFF0;
    // rom_array[3577] = 32'hFFFFFFF1;
    // rom_array[3578] = 32'hFFFFFFF0;
    // rom_array[3579] = 32'hFFFFFFF1;
    // rom_array[3580] = 32'hFFFFFFF0;
    // rom_array[3581] = 32'h000021d9;
    // rom_array[3582] = 32'hFFFFFFF0;
    // rom_array[3583] = 32'h000021e1;
    // rom_array[3584] = 32'hFFFFFFF0;
    // rom_array[3585] = 32'hFFFFFFF1;
    // rom_array[3586] = 32'hFFFFFFF0;
    // rom_array[3587] = 32'hFFFFFFF1;
    // rom_array[3588] = 32'hFFFFFFF0;
    // rom_array[3589] = 32'h000021e9;
    // rom_array[3590] = 32'hFFFFFFF0;
    // rom_array[3591] = 32'h000021f1;
    // rom_array[3592] = 32'hFFFFFFF0;
    // rom_array[3593] = 32'hFFFFFFF1;
    // rom_array[3594] = 32'hFFFFFFF0;
    // rom_array[3595] = 32'hFFFFFFF1;
    // rom_array[3596] = 32'hFFFFFFF0;
    // rom_array[3597] = 32'hFFFFFFF1;
    // rom_array[3598] = 32'hFFFFFFF0;
    // rom_array[3599] = 32'hFFFFFFF1;
    // rom_array[3600] = 32'hFFFFFFF0;
    // rom_array[3601] = 32'hFFFFFFF1;
    // rom_array[3602] = 32'hFFFFFFF0;
    // rom_array[3603] = 32'hFFFFFFF1;
    // rom_array[3604] = 32'hFFFFFFF0;
    // rom_array[3605] = 32'hFFFFFFF1;
    // rom_array[3606] = 32'hFFFFFFF0;
    // rom_array[3607] = 32'hFFFFFFF1;
    // rom_array[3608] = 32'hFFFFFFF0;
    // rom_array[3609] = 32'hFFFFFFF1;
    // rom_array[3610] = 32'hFFFFFFF0;
    // rom_array[3611] = 32'h000021f9;
    // rom_array[3612] = 32'hFFFFFFF0;
    // rom_array[3613] = 32'h00002201;
    // rom_array[3614] = 32'hFFFFFFF0;
    // rom_array[3615] = 32'h00002209;
    // rom_array[3616] = 32'hFFFFFFF0;
    // rom_array[3617] = 32'hFFFFFFF1;
    // rom_array[3618] = 32'hFFFFFFF0;
    // rom_array[3619] = 32'h00002211;
    // rom_array[3620] = 32'hFFFFFFF0;
    // rom_array[3621] = 32'hFFFFFFF1;
    // rom_array[3622] = 32'hFFFFFFF0;
    // rom_array[3623] = 32'h00002219;
    // rom_array[3624] = 32'hFFFFFFF0;
    // rom_array[3625] = 32'h00002221;
    // rom_array[3626] = 32'hFFFFFFF0;
    // rom_array[3627] = 32'h00002229;
    // rom_array[3628] = 32'hFFFFFFF0;
    // rom_array[3629] = 32'h00002231;
    // rom_array[3630] = 32'hFFFFFFF0;
    // rom_array[3631] = 32'h00002239;
    // rom_array[3632] = 32'hFFFFFFF0;
    // rom_array[3633] = 32'h00002241;
    // rom_array[3634] = 32'hFFFFFFF0;
    // rom_array[3635] = 32'h00002249;
    // rom_array[3636] = 32'hFFFFFFF0;
    // rom_array[3637] = 32'h00002251;
    // rom_array[3638] = 32'hFFFFFFF0;
    // rom_array[3639] = 32'h00002259;
    // rom_array[3640] = 32'hFFFFFFF0;
    // rom_array[3641] = 32'hFFFFFFF1;
    // rom_array[3642] = 32'hFFFFFFF0;
    // rom_array[3643] = 32'hFFFFFFF1;
    // rom_array[3644] = 32'hFFFFFFF0;
    // rom_array[3645] = 32'hFFFFFFF1;
    // rom_array[3646] = 32'hFFFFFFF0;
    // rom_array[3647] = 32'hFFFFFFF1;
    // rom_array[3648] = 32'hFFFFFFF0;
    // rom_array[3649] = 32'hFFFFFFF1;
    // rom_array[3650] = 32'hFFFFFFF0;
    // rom_array[3651] = 32'hFFFFFFF1;
    // rom_array[3652] = 32'hFFFFFFF0;
    // rom_array[3653] = 32'hFFFFFFF1;
    // rom_array[3654] = 32'hFFFFFFF0;
    // rom_array[3655] = 32'hFFFFFFF1;
    // rom_array[3656] = 32'hFFFFFFF0;
    // rom_array[3657] = 32'h00002261;
    // rom_array[3658] = 32'hFFFFFFF0;
    // rom_array[3659] = 32'h00002269;
    // rom_array[3660] = 32'hFFFFFFF0;
    // rom_array[3661] = 32'h00002271;
    // rom_array[3662] = 32'hFFFFFFF0;
    // rom_array[3663] = 32'h00002279;
    // rom_array[3664] = 32'hFFFFFFF0;
    // rom_array[3665] = 32'hFFFFFFF1;
    // rom_array[3666] = 32'hFFFFFFF0;
    // rom_array[3667] = 32'h00002281;
    // rom_array[3668] = 32'hFFFFFFF0;
    // rom_array[3669] = 32'hFFFFFFF1;
    // rom_array[3670] = 32'hFFFFFFF0;
    // rom_array[3671] = 32'h00002289;
    // rom_array[3672] = 32'hFFFFFFF0;
    // rom_array[3673] = 32'h00002291;
    // rom_array[3674] = 32'hFFFFFFF0;
    // rom_array[3675] = 32'h00002299;
    // rom_array[3676] = 32'hFFFFFFF0;
    // rom_array[3677] = 32'h000022a1;
    // rom_array[3678] = 32'hFFFFFFF0;
    // rom_array[3679] = 32'h000022a9;
    // rom_array[3680] = 32'hFFFFFFF0;
    // rom_array[3681] = 32'h000022b1;
    // rom_array[3682] = 32'hFFFFFFF0;
    // rom_array[3683] = 32'h000022b9;
    // rom_array[3684] = 32'hFFFFFFF0;
    // rom_array[3685] = 32'h000022c1;
    // rom_array[3686] = 32'hFFFFFFF0;
    // rom_array[3687] = 32'h000022c9;
    // rom_array[3688] = 32'hFFFFFFF0;
    // rom_array[3689] = 32'h000022d1;
    // rom_array[3690] = 32'hFFFFFFF0;
    // rom_array[3691] = 32'h000022d9;
    // rom_array[3692] = 32'hFFFFFFF0;
    // rom_array[3693] = 32'hFFFFFFF0;
    // rom_array[3694] = 32'hFFFFFFF0;
    // rom_array[3695] = 32'hFFFFFFF0;
    // rom_array[3696] = 32'hFFFFFFF0;
    // rom_array[3697] = 32'h000022e1;
    // rom_array[3698] = 32'hFFFFFFF0;
    // rom_array[3699] = 32'h000022e9;
    // rom_array[3700] = 32'hFFFFFFF0;
    // rom_array[3701] = 32'hFFFFFFF0;
    // rom_array[3702] = 32'hFFFFFFF0;
    // rom_array[3703] = 32'hFFFFFFF0;
    // rom_array[3704] = 32'hFFFFFFF0;
    // rom_array[3705] = 32'h000022f1;
    // rom_array[3706] = 32'hFFFFFFF0;
    // rom_array[3707] = 32'h000022f9;
    // rom_array[3708] = 32'hFFFFFFF0;
    // rom_array[3709] = 32'h00002301;
    // rom_array[3710] = 32'hFFFFFFF0;
    // rom_array[3711] = 32'h00002309;
    // rom_array[3712] = 32'hFFFFFFF0;
    // rom_array[3713] = 32'h00002311;
    // rom_array[3714] = 32'hFFFFFFF0;
    // rom_array[3715] = 32'h00002319;
    // rom_array[3716] = 32'hFFFFFFF0;
    // rom_array[3717] = 32'hFFFFFFF0;
    // rom_array[3718] = 32'hFFFFFFF0;
    // rom_array[3719] = 32'hFFFFFFF0;
    // rom_array[3720] = 32'hFFFFFFF0;
    // rom_array[3721] = 32'h00002321;
    // rom_array[3722] = 32'hFFFFFFF0;
    // rom_array[3723] = 32'h00002329;
    // rom_array[3724] = 32'hFFFFFFF0;
    // rom_array[3725] = 32'hFFFFFFF1;
    // rom_array[3726] = 32'hFFFFFFF0;
    // rom_array[3727] = 32'hFFFFFFF1;
    // rom_array[3728] = 32'hFFFFFFF0;
    // rom_array[3729] = 32'h00002331;
    // rom_array[3730] = 32'hFFFFFFF0;
    // rom_array[3731] = 32'h00002339;
    // rom_array[3732] = 32'hFFFFFFF0;
    // rom_array[3733] = 32'hFFFFFFF1;
    // rom_array[3734] = 32'hFFFFFFF0;
    // rom_array[3735] = 32'hFFFFFFF1;
    // rom_array[3736] = 32'hFFFFFFF0;
    // rom_array[3737] = 32'h00002341;
    // rom_array[3738] = 32'hFFFFFFF0;
    // rom_array[3739] = 32'h00002349;
    // rom_array[3740] = 32'hFFFFFFF0;
    // rom_array[3741] = 32'h00002351;
    // rom_array[3742] = 32'hFFFFFFF0;
    // rom_array[3743] = 32'hFFFFFFF0;
    // rom_array[3744] = 32'hFFFFFFF0;
    // rom_array[3745] = 32'h00002359;
    // rom_array[3746] = 32'hFFFFFFF0;
    // rom_array[3747] = 32'h00002361;
    // rom_array[3748] = 32'hFFFFFFF0;
    // rom_array[3749] = 32'hFFFFFFF0;
    // rom_array[3750] = 32'hFFFFFFF0;
    // rom_array[3751] = 32'h00002369;
    // rom_array[3752] = 32'hFFFFFFF0;
    // rom_array[3753] = 32'h00002371;
    // rom_array[3754] = 32'hFFFFFFF0;
    // rom_array[3755] = 32'h00002379;
    // rom_array[3756] = 32'hFFFFFFF0;
    // rom_array[3757] = 32'hFFFFFFF1;
    // rom_array[3758] = 32'hFFFFFFF0;
    // rom_array[3759] = 32'h00002381;
    // rom_array[3760] = 32'hFFFFFFF0;
    // rom_array[3761] = 32'h00002389;
    // rom_array[3762] = 32'hFFFFFFF0;
    // rom_array[3763] = 32'h00002391;
    // rom_array[3764] = 32'hFFFFFFF0;
    // rom_array[3765] = 32'hFFFFFFF1;
    // rom_array[3766] = 32'hFFFFFFF0;
    // rom_array[3767] = 32'h00002399;
    // rom_array[3768] = 32'hFFFFFFF0;
    // rom_array[3769] = 32'h000023a1;
    // rom_array[3770] = 32'hFFFFFFF0;
    // rom_array[3771] = 32'hFFFFFFF0;
    // rom_array[3772] = 32'hFFFFFFF0;
    // rom_array[3773] = 32'h000023a9;
    // rom_array[3774] = 32'hFFFFFFF0;
    // rom_array[3775] = 32'h000023b1;
    // rom_array[3776] = 32'hFFFFFFF0;
    // rom_array[3777] = 32'hFFFFFFF0;
    // rom_array[3778] = 32'hFFFFFFF0;
    // rom_array[3779] = 32'h000023b9;
    // rom_array[3780] = 32'hFFFFFFF0;
    // rom_array[3781] = 32'h000023c1;
    // rom_array[3782] = 32'hFFFFFFF0;
    // rom_array[3783] = 32'h000023c9;
    // rom_array[3784] = 32'hFFFFFFF0;
    // rom_array[3785] = 32'h000023d1;
    // rom_array[3786] = 32'hFFFFFFF0;
    // rom_array[3787] = 32'hFFFFFFF1;
    // rom_array[3788] = 32'hFFFFFFF0;
    // rom_array[3789] = 32'h000023d9;
    // rom_array[3790] = 32'hFFFFFFF0;
    // rom_array[3791] = 32'h000023e1;
    // rom_array[3792] = 32'hFFFFFFF0;
    // rom_array[3793] = 32'hFFFFFFF1;
    // rom_array[3794] = 32'hFFFFFFF0;
    // rom_array[3795] = 32'h000023e9;
    // rom_array[3796] = 32'hFFFFFFF0;
    // rom_array[3797] = 32'h000023f1;
    // rom_array[3798] = 32'hFFFFFFF0;
    // rom_array[3799] = 32'h000023f9;
    // rom_array[3800] = 32'hFFFFFFF0;
    // rom_array[3801] = 32'hFFFFFFF1;
    // rom_array[3802] = 32'hFFFFFFF0;
    // rom_array[3803] = 32'h00002401;
    // rom_array[3804] = 32'hFFFFFFF0;
    // rom_array[3805] = 32'hFFFFFFF1;
    // rom_array[3806] = 32'hFFFFFFF0;
    // rom_array[3807] = 32'h00002409;
    // rom_array[3808] = 32'hFFFFFFF0;
    // rom_array[3809] = 32'h00002411;
    // rom_array[3810] = 32'hFFFFFFF0;
    // rom_array[3811] = 32'h00002419;
    // rom_array[3812] = 32'hFFFFFFF0;
    // rom_array[3813] = 32'hFFFFFFF0;
    // rom_array[3814] = 32'hFFFFFFF0;
    // rom_array[3815] = 32'hFFFFFFF0;
    // rom_array[3816] = 32'hFFFFFFF0;
    // rom_array[3817] = 32'hFFFFFFF0;
    // rom_array[3818] = 32'hFFFFFFF0;
    // rom_array[3819] = 32'hFFFFFFF0;
    // rom_array[3820] = 32'hFFFFFFF0;
    // rom_array[3821] = 32'h00002421;
    // rom_array[3822] = 32'hFFFFFFF0;
    // rom_array[3823] = 32'h00002429;
    // rom_array[3824] = 32'hFFFFFFF0;
    // rom_array[3825] = 32'hFFFFFFF0;
    // rom_array[3826] = 32'hFFFFFFF0;
    // rom_array[3827] = 32'hFFFFFFF0;
    // rom_array[3828] = 32'hFFFFFFF0;
    // rom_array[3829] = 32'h00002431;
    // rom_array[3830] = 32'hFFFFFFF0;
    // rom_array[3831] = 32'h00002439;
    // rom_array[3832] = 32'hFFFFFFF0;
    // rom_array[3833] = 32'hFFFFFFF1;
    // rom_array[3834] = 32'hFFFFFFF0;
    // rom_array[3835] = 32'hFFFFFFF1;
    // rom_array[3836] = 32'hFFFFFFF0;
    // rom_array[3837] = 32'h00002441;
    // rom_array[3838] = 32'hFFFFFFF0;
    // rom_array[3839] = 32'h00002449;
    // rom_array[3840] = 32'hFFFFFFF0;
    // rom_array[3841] = 32'hFFFFFFF1;
    // rom_array[3842] = 32'hFFFFFFF0;
    // rom_array[3843] = 32'hFFFFFFF1;
    // rom_array[3844] = 32'hFFFFFFF0;
    // rom_array[3845] = 32'h00002451;
    // rom_array[3846] = 32'hFFFFFFF0;
    // rom_array[3847] = 32'h00002459;
    // rom_array[3848] = 32'hFFFFFFF0;
    // rom_array[3849] = 32'hFFFFFFF0;
    // rom_array[3850] = 32'hFFFFFFF0;
    // rom_array[3851] = 32'hFFFFFFF0;
    // rom_array[3852] = 32'hFFFFFFF0;
    // rom_array[3853] = 32'h00002461;
    // rom_array[3854] = 32'hFFFFFFF0;
    // rom_array[3855] = 32'h00002469;
    // rom_array[3856] = 32'hFFFFFFF0;
    // rom_array[3857] = 32'hFFFFFFF1;
    // rom_array[3858] = 32'hFFFFFFF0;
    // rom_array[3859] = 32'h00002471;
    // rom_array[3860] = 32'hFFFFFFF0;
    // rom_array[3861] = 32'h00002479;
    // rom_array[3862] = 32'hFFFFFFF0;
    // rom_array[3863] = 32'h00002481;
    // rom_array[3864] = 32'hFFFFFFF0;
    // rom_array[3865] = 32'h00002489;
    // rom_array[3866] = 32'hFFFFFFF0;
    // rom_array[3867] = 32'hFFFFFFF0;
    // rom_array[3868] = 32'hFFFFFFF0;
    // rom_array[3869] = 32'h00002491;
    // rom_array[3870] = 32'hFFFFFFF0;
    // rom_array[3871] = 32'hFFFFFFF0;
    // rom_array[3872] = 32'hFFFFFFF0;
    // rom_array[3873] = 32'hFFFFFFF0;
    // rom_array[3874] = 32'hFFFFFFF0;
    // rom_array[3875] = 32'h00002499;
    // rom_array[3876] = 32'hFFFFFFF0;
    // rom_array[3877] = 32'hFFFFFFF0;
    // rom_array[3878] = 32'hFFFFFFF0;
    // rom_array[3879] = 32'h000024a1;
    // rom_array[3880] = 32'hFFFFFFF0;
    // rom_array[3881] = 32'h000024a9;
    // rom_array[3882] = 32'hFFFFFFF0;
    // rom_array[3883] = 32'hFFFFFFF0;
    // rom_array[3884] = 32'hFFFFFFF0;
    // rom_array[3885] = 32'h000024b1;
    // rom_array[3886] = 32'hFFFFFFF0;
    // rom_array[3887] = 32'hFFFFFFF0;
    // rom_array[3888] = 32'hFFFFFFF0;
    // rom_array[3889] = 32'hFFFFFFF0;
    // rom_array[3890] = 32'hFFFFFFF0;
    // rom_array[3891] = 32'h000024b9;
    // rom_array[3892] = 32'hFFFFFFF0;
    // rom_array[3893] = 32'hFFFFFFF0;
    // rom_array[3894] = 32'hFFFFFFF0;
    // rom_array[3895] = 32'h000024c1;
    // rom_array[3896] = 32'hFFFFFFF0;
    // rom_array[3897] = 32'hFFFFFFF1;
    // rom_array[3898] = 32'hFFFFFFF0;
    // rom_array[3899] = 32'h000024c9;
    // rom_array[3900] = 32'hFFFFFFF0;
    // rom_array[3901] = 32'hFFFFFFF1;
    // rom_array[3902] = 32'hFFFFFFF0;
    // rom_array[3903] = 32'h000024d1;
    // rom_array[3904] = 32'hFFFFFFF0;
    // rom_array[3905] = 32'hFFFFFFF1;
    // rom_array[3906] = 32'hFFFFFFF0;
    // rom_array[3907] = 32'h000024d9;
    // rom_array[3908] = 32'hFFFFFFF0;
    // rom_array[3909] = 32'hFFFFFFF1;
    // rom_array[3910] = 32'hFFFFFFF0;
    // rom_array[3911] = 32'h000024e1;
    // rom_array[3912] = 32'hFFFFFFF0;
    // rom_array[3913] = 32'hFFFFFFF0;
    // rom_array[3914] = 32'h000024e9;
    // rom_array[3915] = 32'hFFFFFFF0;
    // rom_array[3916] = 32'h000024f1;
    // rom_array[3917] = 32'hFFFFFFF0;
    // rom_array[3918] = 32'hFFFFFFF0;
    // rom_array[3919] = 32'hFFFFFFF0;
    // rom_array[3920] = 32'hFFFFFFF0;
    // rom_array[3921] = 32'hFFFFFFF0;
    // rom_array[3922] = 32'h000024f9;
    // rom_array[3923] = 32'hFFFFFFF0;
    // rom_array[3924] = 32'hFFFFFFF0;
    // rom_array[3925] = 32'hFFFFFFF0;
    // rom_array[3926] = 32'hFFFFFFF0;
    // rom_array[3927] = 32'hFFFFFFF0;
    // rom_array[3928] = 32'hFFFFFFF0;
    // rom_array[3929] = 32'hFFFFFFF0;
    // rom_array[3930] = 32'h00002501;
    // rom_array[3931] = 32'hFFFFFFF0;
    // rom_array[3932] = 32'h00002509;
    // rom_array[3933] = 32'hFFFFFFF0;
    // rom_array[3934] = 32'hFFFFFFF0;
    // rom_array[3935] = 32'hFFFFFFF0;
    // rom_array[3936] = 32'hFFFFFFF0;
    // rom_array[3937] = 32'hFFFFFFF0;
    // rom_array[3938] = 32'hFFFFFFF0;
    // rom_array[3939] = 32'hFFFFFFF0;
    // rom_array[3940] = 32'hFFFFFFF0;
    // rom_array[3941] = 32'hFFFFFFF0;
    // rom_array[3942] = 32'h00002511;
    // rom_array[3943] = 32'hFFFFFFF0;
    // rom_array[3944] = 32'h00002519;
    // rom_array[3945] = 32'hFFFFFFF0;
    // rom_array[3946] = 32'h00002521;
    // rom_array[3947] = 32'hFFFFFFF0;
    // rom_array[3948] = 32'hFFFFFFF1;
    // rom_array[3949] = 32'hFFFFFFF0;
    // rom_array[3950] = 32'h00002529;
    // rom_array[3951] = 32'hFFFFFFF0;
    // rom_array[3952] = 32'h00002531;
    // rom_array[3953] = 32'hFFFFFFF0;
    // rom_array[3954] = 32'hFFFFFFF0;
    // rom_array[3955] = 32'hFFFFFFF0;
    // rom_array[3956] = 32'hFFFFFFF0;
    // rom_array[3957] = 32'hFFFFFFF0;
    // rom_array[3958] = 32'h00002539;
    // rom_array[3959] = 32'hFFFFFFF0;
    // rom_array[3960] = 32'h00002541;
    // rom_array[3961] = 32'hFFFFFFF0;
    // rom_array[3962] = 32'hFFFFFFF0;
    // rom_array[3963] = 32'hFFFFFFF0;
    // rom_array[3964] = 32'hFFFFFFF0;
    // rom_array[3965] = 32'hFFFFFFF0;
    // rom_array[3966] = 32'h00002549;
    // rom_array[3967] = 32'hFFFFFFF0;
    // rom_array[3968] = 32'h00002551;
    // rom_array[3969] = 32'hFFFFFFF0;
    // rom_array[3970] = 32'hFFFFFFF1;
    // rom_array[3971] = 32'hFFFFFFF0;
    // rom_array[3972] = 32'hFFFFFFF1;
    // rom_array[3973] = 32'hFFFFFFF0;
    // rom_array[3974] = 32'h00002559;
    // rom_array[3975] = 32'hFFFFFFF0;
    // rom_array[3976] = 32'h00002561;
    // rom_array[3977] = 32'hFFFFFFF0;
    // rom_array[3978] = 32'hFFFFFFF1;
    // rom_array[3979] = 32'hFFFFFFF0;
    // rom_array[3980] = 32'hFFFFFFF1;
    // rom_array[3981] = 32'hFFFFFFF0;
    // rom_array[3982] = 32'h00002569;
    // rom_array[3983] = 32'hFFFFFFF0;
    // rom_array[3984] = 32'h00002571;
    // rom_array[3985] = 32'hFFFFFFF0;
    // rom_array[3986] = 32'hFFFFFFF0;
    // rom_array[3987] = 32'hFFFFFFF0;
    // rom_array[3988] = 32'hFFFFFFF0;
    // rom_array[3989] = 32'hFFFFFFF0;
    // rom_array[3990] = 32'h00002579;
    // rom_array[3991] = 32'hFFFFFFF0;
    // rom_array[3992] = 32'h00002581;
    // rom_array[3993] = 32'hFFFFFFF0;
    // rom_array[3994] = 32'h00002589;
    // rom_array[3995] = 32'hFFFFFFF0;
    // rom_array[3996] = 32'h00002591;
    // rom_array[3997] = 32'hFFFFFFF0;
    // rom_array[3998] = 32'h00002599;
    // rom_array[3999] = 32'hFFFFFFF0;
    // rom_array[4000] = 32'h000025a1;
    // rom_array[4001] = 32'hFFFFFFF0;
    // rom_array[4002] = 32'hFFFFFFF0;
    // rom_array[4003] = 32'hFFFFFFF0;
    // rom_array[4004] = 32'hFFFFFFF0;
    // rom_array[4005] = 32'hFFFFFFF0;
    // rom_array[4006] = 32'h000025a9;
    // rom_array[4007] = 32'hFFFFFFF0;
    // rom_array[4008] = 32'h000025b1;
    // rom_array[4009] = 32'hFFFFFFF0;
    // rom_array[4010] = 32'h000025b9;
    // rom_array[4011] = 32'hFFFFFFF0;
    // rom_array[4012] = 32'hFFFFFFF1;
    // rom_array[4013] = 32'hFFFFFFF0;
    // rom_array[4014] = 32'h000025c1;
    // rom_array[4015] = 32'hFFFFFFF0;
    // rom_array[4016] = 32'h000025c9;
    // rom_array[4017] = 32'hFFFFFFF0;
    // rom_array[4018] = 32'hFFFFFFF1;
    // rom_array[4019] = 32'hFFFFFFF0;
    // rom_array[4020] = 32'hFFFFFFF1;
    // rom_array[4021] = 32'hFFFFFFF0;
    // rom_array[4022] = 32'hFFFFFFF1;
    // rom_array[4023] = 32'hFFFFFFF0;
    // rom_array[4024] = 32'hFFFFFFF1;
    // rom_array[4025] = 32'hFFFFFFF0;
    // rom_array[4026] = 32'h000025d1;
    // rom_array[4027] = 32'hFFFFFFF0;
    // rom_array[4028] = 32'h000025d9;
    // rom_array[4029] = 32'hFFFFFFF0;
    // rom_array[4030] = 32'h000025e1;
    // rom_array[4031] = 32'hFFFFFFF0;
    // rom_array[4032] = 32'h000025e9;
    // rom_array[4033] = 32'hFFFFFFF0;
    // rom_array[4034] = 32'h000025f1;
    // rom_array[4035] = 32'hFFFFFFF0;
    // rom_array[4036] = 32'h000025f9;
    // rom_array[4037] = 32'hFFFFFFF0;
    // rom_array[4038] = 32'hFFFFFFF0;
    // rom_array[4039] = 32'hFFFFFFF0;
    // rom_array[4040] = 32'hFFFFFFF0;
    // rom_array[4041] = 32'hFFFFFFF0;
    // rom_array[4042] = 32'h00002601;
    // rom_array[4043] = 32'hFFFFFFF0;
    // rom_array[4044] = 32'h00002609;
    // rom_array[4045] = 32'hFFFFFFF0;
    // rom_array[4046] = 32'hFFFFFFF0;
    // rom_array[4047] = 32'hFFFFFFF0;
    // rom_array[4048] = 32'hFFFFFFF0;
    // rom_array[4049] = 32'hFFFFFFF0;
    // rom_array[4050] = 32'h00002611;
    // rom_array[4051] = 32'hFFFFFFF0;
    // rom_array[4052] = 32'h00002619;
    // rom_array[4053] = 32'hFFFFFFF0;
    // rom_array[4054] = 32'hFFFFFFF0;
    // rom_array[4055] = 32'hFFFFFFF0;
    // rom_array[4056] = 32'hFFFFFFF0;
    // rom_array[4057] = 32'hFFFFFFF0;
    // rom_array[4058] = 32'h00002621;
    // rom_array[4059] = 32'hFFFFFFF0;
    // rom_array[4060] = 32'h00002629;
    // rom_array[4061] = 32'hFFFFFFF0;
    // rom_array[4062] = 32'h00002631;
    // rom_array[4063] = 32'hFFFFFFF0;
    // rom_array[4064] = 32'hFFFFFFF1;
    // rom_array[4065] = 32'hFFFFFFF0;
    // rom_array[4066] = 32'h00002639;
    // rom_array[4067] = 32'hFFFFFFF0;
    // rom_array[4068] = 32'hFFFFFFF1;
    // rom_array[4069] = 32'hFFFFFFF0;
    // rom_array[4070] = 32'h00002641;
    // rom_array[4071] = 32'hFFFFFFF0;
    // rom_array[4072] = 32'hFFFFFFF1;
    // rom_array[4073] = 32'hFFFFFFF0;
    // rom_array[4074] = 32'h00002649;
    // rom_array[4075] = 32'hFFFFFFF0;
    // rom_array[4076] = 32'hFFFFFFF0;
    // rom_array[4077] = 32'hFFFFFFF0;
    // rom_array[4078] = 32'h00002651;
    // rom_array[4079] = 32'hFFFFFFF0;
    // rom_array[4080] = 32'hFFFFFFF0;
    // rom_array[4081] = 32'hFFFFFFF0;
    // rom_array[4082] = 32'h00002659;
    // rom_array[4083] = 32'hFFFFFFF0;
    // rom_array[4084] = 32'hFFFFFFF0;
    // rom_array[4085] = 32'hFFFFFFF0;
    // rom_array[4086] = 32'h00002661;
    // rom_array[4087] = 32'hFFFFFFF0;
    // rom_array[4088] = 32'h00002669;
    // rom_array[4089] = 32'hFFFFFFF0;
    // rom_array[4090] = 32'hFFFFFFF0;
    // rom_array[4091] = 32'hFFFFFFF0;
    // rom_array[4092] = 32'hFFFFFFF0;
    // rom_array[4093] = 32'hFFFFFFF0;
    // rom_array[4094] = 32'h00002671;
    // rom_array[4095] = 32'hFFFFFFF0;
    // rom_array[4096] = 32'h00002679;
    // rom_array[4097] = 32'hFFFFFFF0;
    // rom_array[4098] = 32'h00002681;
    // rom_array[4099] = 32'hFFFFFFF0;
    // rom_array[4100] = 32'hFFFFFFF1;
    // rom_array[4101] = 32'hFFFFFFF0;
    // rom_array[4102] = 32'h00002689;
    // rom_array[4103] = 32'hFFFFFFF0;
    // rom_array[4104] = 32'hFFFFFFF1;
    // rom_array[4105] = 32'hFFFFFFF0;
    // rom_array[4106] = 32'h00002691;
    // rom_array[4107] = 32'hFFFFFFF0;
    // rom_array[4108] = 32'hFFFFFFF1;
    // rom_array[4109] = 32'hFFFFFFF0;
    // rom_array[4110] = 32'h00002699;
    // rom_array[4111] = 32'hFFFFFFF0;
    // rom_array[4112] = 32'h000026a1;
    // rom_array[4113] = 32'hFFFFFFF0;
    // rom_array[4114] = 32'h000026a9;
    // rom_array[4115] = 32'hFFFFFFF0;
    // rom_array[4116] = 32'hFFFFFFF1;
    // rom_array[4117] = 32'hFFFFFFF0;
    // rom_array[4118] = 32'h000026b1;
    // rom_array[4119] = 32'hFFFFFFF0;
    // rom_array[4120] = 32'h000026b9;
    // rom_array[4121] = 32'hFFFFFFF0;
    // rom_array[4122] = 32'hFFFFFFF1;
    // rom_array[4123] = 32'hFFFFFFF0;
    // rom_array[4124] = 32'hFFFFFFF1;
    // rom_array[4125] = 32'hFFFFFFF0;
    // rom_array[4126] = 32'h000026c1;
    // rom_array[4127] = 32'hFFFFFFF0;
    // rom_array[4128] = 32'h000026c9;
    // rom_array[4129] = 32'hFFFFFFF0;
    // rom_array[4130] = 32'h000026d1;
    // rom_array[4131] = 32'hFFFFFFF0;
    // rom_array[4132] = 32'hFFFFFFF0;
    // rom_array[4133] = 32'hFFFFFFF0;
    // rom_array[4134] = 32'h000026d9;
    // rom_array[4135] = 32'hFFFFFFF0;
    // rom_array[4136] = 32'hFFFFFFF0;
    // rom_array[4137] = 32'hFFFFFFF0;
    // rom_array[4138] = 32'h000026e1;
    // rom_array[4139] = 32'hFFFFFFF0;
    // rom_array[4140] = 32'h000026e9;
    // rom_array[4141] = 32'hFFFFFFF0;
    // rom_array[4142] = 32'h000026f1;
    // rom_array[4143] = 32'hFFFFFFF0;
    // rom_array[4144] = 32'h000026f9;
    // rom_array[4145] = 32'hFFFFFFF0;
    // rom_array[4146] = 32'h00002701;
    // rom_array[4147] = 32'hFFFFFFF0;
    // rom_array[4148] = 32'h00002709;
    // rom_array[4149] = 32'hFFFFFFF0;
    // rom_array[4150] = 32'h00002711;
    // rom_array[4151] = 32'hFFFFFFF0;
    // rom_array[4152] = 32'hFFFFFFF1;
    // rom_array[4153] = 32'hFFFFFFF0;
    // rom_array[4154] = 32'h00002719;
    // rom_array[4155] = 32'hFFFFFFF0;
    // rom_array[4156] = 32'h00002721;
    // rom_array[4157] = 32'hFFFFFFF0;
    // rom_array[4158] = 32'hFFFFFFF1;
    // rom_array[4159] = 32'hFFFFFFF0;
    // rom_array[4160] = 32'hFFFFFFF1;
    // rom_array[4161] = 32'hFFFFFFF0;
    // rom_array[4162] = 32'h00002729;
    // rom_array[4163] = 32'hFFFFFFF0;
    // rom_array[4164] = 32'h00002731;
    // rom_array[4165] = 32'hFFFFFFF0;
    // rom_array[4166] = 32'hFFFFFFF1;
    // rom_array[4167] = 32'hFFFFFFF0;
    // rom_array[4168] = 32'hFFFFFFF1;
    // rom_array[4169] = 32'hFFFFFFF0;
    // rom_array[4170] = 32'h00002739;
    // rom_array[4171] = 32'hFFFFFFF0;
    // rom_array[4172] = 32'h00002741;
    // rom_array[4173] = 32'hFFFFFFF0;
    // rom_array[4174] = 32'h00002749;
    // rom_array[4175] = 32'hFFFFFFF0;
    // rom_array[4176] = 32'hFFFFFFF1;
    // rom_array[4177] = 32'hFFFFFFF0;
    // rom_array[4178] = 32'h00002751;
    // rom_array[4179] = 32'hFFFFFFF0;
    // rom_array[4180] = 32'hFFFFFFF1;
    // rom_array[4181] = 32'hFFFFFFF0;
    // rom_array[4182] = 32'h00002759;
    // rom_array[4183] = 32'hFFFFFFF0;
    // rom_array[4184] = 32'hFFFFFFF1;
    // rom_array[4185] = 32'hFFFFFFF0;
    // rom_array[4186] = 32'h00002761;
    // rom_array[4187] = 32'hFFFFFFF0;
    // rom_array[4188] = 32'h00002769;
    // rom_array[4189] = 32'hFFFFFFF0;
    // rom_array[4190] = 32'h00002771;
    // rom_array[4191] = 32'hFFFFFFF0;
    // rom_array[4192] = 32'hFFFFFFF1;
    // rom_array[4193] = 32'hFFFFFFF0;
    // rom_array[4194] = 32'h00002779;
    // rom_array[4195] = 32'hFFFFFFF0;
    // rom_array[4196] = 32'h00002781;
    // rom_array[4197] = 32'hFFFFFFF0;
    // rom_array[4198] = 32'h00002789;
    // rom_array[4199] = 32'hFFFFFFF0;
    // rom_array[4200] = 32'hFFFFFFF1;
    // rom_array[4201] = 32'hFFFFFFF0;
    // rom_array[4202] = 32'h00002791;
    // rom_array[4203] = 32'hFFFFFFF0;
    // rom_array[4204] = 32'h00002799;
    // rom_array[4205] = 32'hFFFFFFF0;
    // rom_array[4206] = 32'h000027a1;
    // rom_array[4207] = 32'hFFFFFFF0;
    // rom_array[4208] = 32'hFFFFFFF1;
    // rom_array[4209] = 32'hFFFFFFF0;
    // rom_array[4210] = 32'h000027a9;
    // rom_array[4211] = 32'hFFFFFFF0;
    // rom_array[4212] = 32'h000027b1;
    // rom_array[4213] = 32'hFFFFFFF0;
    // rom_array[4214] = 32'h000027b9;
    // rom_array[4215] = 32'hFFFFFFF0;
    // rom_array[4216] = 32'hFFFFFFF1;
    // rom_array[4217] = 32'hFFFFFFF0;
    // rom_array[4218] = 32'h000027c1;
    // rom_array[4219] = 32'hFFFFFFF0;
    // rom_array[4220] = 32'h000027c9;
    // rom_array[4221] = 32'hFFFFFFF0;
    // rom_array[4222] = 32'h000027d1;
    // rom_array[4223] = 32'hFFFFFFF0;
    // rom_array[4224] = 32'h000027d9;
    // rom_array[4225] = 32'hFFFFFFF0;
    // rom_array[4226] = 32'h000027e1;
    // rom_array[4227] = 32'hFFFFFFF0;
    // rom_array[4228] = 32'h000027e9;
    // rom_array[4229] = 32'hFFFFFFF0;
    // rom_array[4230] = 32'h000027f1;
    // rom_array[4231] = 32'hFFFFFFF0;
    // rom_array[4232] = 32'hFFFFFFF1;
    // rom_array[4233] = 32'hFFFFFFF0;
    // rom_array[4234] = 32'h000027f9;
    // rom_array[4235] = 32'hFFFFFFF0;
    // rom_array[4236] = 32'h00002801;
    // rom_array[4237] = 32'hFFFFFFF0;
    // rom_array[4238] = 32'h00002809;
    // rom_array[4239] = 32'hFFFFFFF0;
    // rom_array[4240] = 32'h00002811;
    // rom_array[4241] = 32'hFFFFFFF0;
    // rom_array[4242] = 32'h00002819;
    // rom_array[4243] = 32'hFFFFFFF0;
    // rom_array[4244] = 32'h00002821;
    // rom_array[4245] = 32'hFFFFFFF0;
    // rom_array[4246] = 32'hFFFFFFF0;
    // rom_array[4247] = 32'hFFFFFFF0;
    // rom_array[4248] = 32'hFFFFFFF0;
    // rom_array[4249] = 32'hFFFFFFF0;
    // rom_array[4250] = 32'hFFFFFFF1;
    // rom_array[4251] = 32'hFFFFFFF0;
    // rom_array[4252] = 32'hFFFFFFF1;
    // rom_array[4253] = 32'hFFFFFFF0;
    // rom_array[4254] = 32'hFFFFFFF1;
    // rom_array[4255] = 32'hFFFFFFF0;
    // rom_array[4256] = 32'hFFFFFFF1;
    // rom_array[4257] = 32'hFFFFFFF0;
    // rom_array[4258] = 32'hFFFFFFF1;
    // rom_array[4259] = 32'hFFFFFFF0;
    // rom_array[4260] = 32'hFFFFFFF1;
    // rom_array[4261] = 32'hFFFFFFF0;
    // rom_array[4262] = 32'hFFFFFFF1;
    // rom_array[4263] = 32'hFFFFFFF0;
    // rom_array[4264] = 32'hFFFFFFF1;
    // rom_array[4265] = 32'hFFFFFFF0;
    // rom_array[4266] = 32'h00002829;
    // rom_array[4267] = 32'hFFFFFFF0;
    // rom_array[4268] = 32'h00002831;
    // rom_array[4269] = 32'hFFFFFFF0;
    // rom_array[4270] = 32'hFFFFFFF0;
    // rom_array[4271] = 32'hFFFFFFF0;
    // rom_array[4272] = 32'hFFFFFFF0;
    // rom_array[4273] = 32'hFFFFFFF0;
    // rom_array[4274] = 32'h00002839;
    // rom_array[4275] = 32'hFFFFFFF0;
    // rom_array[4276] = 32'h00002841;
    // rom_array[4277] = 32'hFFFFFFF0;
    // rom_array[4278] = 32'hFFFFFFF0;
    // rom_array[4279] = 32'hFFFFFFF0;
    // rom_array[4280] = 32'hFFFFFFF0;
    // rom_array[4281] = 32'hFFFFFFF0;
    // rom_array[4282] = 32'h00002849;
    // rom_array[4283] = 32'hFFFFFFF0;
    // rom_array[4284] = 32'h00002851;
    // rom_array[4285] = 32'hFFFFFFF0;
    // rom_array[4286] = 32'h00002859;
    // rom_array[4287] = 32'hFFFFFFF0;
    // rom_array[4288] = 32'hFFFFFFF1;
    // rom_array[4289] = 32'hFFFFFFF0;
    // rom_array[4290] = 32'h00002861;
    // rom_array[4291] = 32'hFFFFFFF0;
    // rom_array[4292] = 32'h00002869;
    // rom_array[4293] = 32'hFFFFFFF0;
    // rom_array[4294] = 32'hFFFFFFF1;
    // rom_array[4295] = 32'hFFFFFFF0;
    // rom_array[4296] = 32'hFFFFFFF1;
    // rom_array[4297] = 32'hFFFFFFF0;
    // rom_array[4298] = 32'h00002871;
    // rom_array[4299] = 32'hFFFFFFF0;
    // rom_array[4300] = 32'h00002879;
    // rom_array[4301] = 32'hFFFFFFF0;
    // rom_array[4302] = 32'hFFFFFFF1;
    // rom_array[4303] = 32'hFFFFFFF0;
    // rom_array[4304] = 32'hFFFFFFF1;
    // rom_array[4305] = 32'hFFFFFFF0;
    // rom_array[4306] = 32'h00002881;
    // rom_array[4307] = 32'hFFFFFFF0;
    // rom_array[4308] = 32'h00002889;
    // rom_array[4309] = 32'hFFFFFFF0;
    // rom_array[4310] = 32'h00002891;
    // rom_array[4311] = 32'hFFFFFFF0;
    // rom_array[4312] = 32'hFFFFFFF1;
    // rom_array[4313] = 32'hFFFFFFF0;
    // rom_array[4314] = 32'h00002899;
    // rom_array[4315] = 32'hFFFFFFF0;
    // rom_array[4316] = 32'hFFFFFFF1;
    // rom_array[4317] = 32'hFFFFFFF0;
    // rom_array[4318] = 32'h000028a1;
    // rom_array[4319] = 32'hFFFFFFF0;
    // rom_array[4320] = 32'hFFFFFFF1;
    // rom_array[4321] = 32'hFFFFFFF0;
    // rom_array[4322] = 32'h000028a9;
    // rom_array[4323] = 32'hFFFFFFF0;
    // rom_array[4324] = 32'h000028b1;
    // rom_array[4325] = 32'hFFFFFFF0;
    // rom_array[4326] = 32'h000028b9;
    // rom_array[4327] = 32'hFFFFFFF0;
    // rom_array[4328] = 32'hFFFFFFF0;
    // rom_array[4329] = 32'hFFFFFFF0;
    // rom_array[4330] = 32'h000028c1;
    // rom_array[4331] = 32'hFFFFFFF0;
    // rom_array[4332] = 32'h000028c9;
    // rom_array[4333] = 32'hFFFFFFF0;
    // rom_array[4334] = 32'hFFFFFFF0;
    // rom_array[4335] = 32'hFFFFFFF0;
    // rom_array[4336] = 32'hFFFFFFF0;
    // rom_array[4337] = 32'hFFFFFFF0;
    // rom_array[4338] = 32'h000028d1;
    // rom_array[4339] = 32'hFFFFFFF0;
    // rom_array[4340] = 32'hFFFFFFF0;
    // rom_array[4341] = 32'hFFFFFFF0;
    // rom_array[4342] = 32'h000028d9;
    // rom_array[4343] = 32'hFFFFFFF0;
    // rom_array[4344] = 32'hFFFFFFF0;
    // rom_array[4345] = 32'hFFFFFFF0;
    // rom_array[4346] = 32'h000028e1;
    // rom_array[4347] = 32'hFFFFFFF0;
    // rom_array[4348] = 32'hFFFFFFF1;
    // rom_array[4349] = 32'hFFFFFFF0;
    // rom_array[4350] = 32'h000028e9;
    // rom_array[4351] = 32'hFFFFFFF0;
    // rom_array[4352] = 32'h000028f1;
    // rom_array[4353] = 32'hFFFFFFF0;
    // rom_array[4354] = 32'h000028f9;
    // rom_array[4355] = 32'hFFFFFFF0;
    // rom_array[4356] = 32'hFFFFFFF0;
    // rom_array[4357] = 32'hFFFFFFF0;
    // rom_array[4358] = 32'h00002901;
    // rom_array[4359] = 32'hFFFFFFF0;
    // rom_array[4360] = 32'hFFFFFFF0;
    // rom_array[4361] = 32'h00002909;
    // rom_array[4362] = 32'hFFFFFFF0;
    // rom_array[4363] = 32'h00002911;
    // rom_array[4364] = 32'hFFFFFFF0;
    // rom_array[4365] = 32'hFFFFFFF0;
    // rom_array[4366] = 32'hFFFFFFF0;
    // rom_array[4367] = 32'hFFFFFFF0;
    // rom_array[4368] = 32'hFFFFFFF0;
    // rom_array[4369] = 32'h00002919;
    // rom_array[4370] = 32'hFFFFFFF0;
    // rom_array[4371] = 32'hFFFFFFF0;
    // rom_array[4372] = 32'hFFFFFFF0;
    // rom_array[4373] = 32'hFFFFFFF0;
    // rom_array[4374] = 32'hFFFFFFF0;
    // rom_array[4375] = 32'hFFFFFFF0;
    // rom_array[4376] = 32'hFFFFFFF0;
    // rom_array[4377] = 32'h00002921;
    // rom_array[4378] = 32'hFFFFFFF0;
    // rom_array[4379] = 32'h00002929;
    // rom_array[4380] = 32'hFFFFFFF0;
    // rom_array[4381] = 32'hFFFFFFF0;
    // rom_array[4382] = 32'hFFFFFFF0;
    // rom_array[4383] = 32'hFFFFFFF0;
    // rom_array[4384] = 32'hFFFFFFF0;
    // rom_array[4385] = 32'hFFFFFFF0;
    // rom_array[4386] = 32'hFFFFFFF0;
    // rom_array[4387] = 32'hFFFFFFF0;
    // rom_array[4388] = 32'hFFFFFFF0;
    // rom_array[4389] = 32'h00002931;
    // rom_array[4390] = 32'hFFFFFFF0;
    // rom_array[4391] = 32'h00002939;
    // rom_array[4392] = 32'hFFFFFFF0;
    // rom_array[4393] = 32'h00002941;
    // rom_array[4394] = 32'hFFFFFFF0;
    // rom_array[4395] = 32'hFFFFFFF1;
    // rom_array[4396] = 32'hFFFFFFF0;
    // rom_array[4397] = 32'h00002949;
    // rom_array[4398] = 32'hFFFFFFF0;
    // rom_array[4399] = 32'h00002951;
    // rom_array[4400] = 32'hFFFFFFF0;
    // rom_array[4401] = 32'hFFFFFFF0;
    // rom_array[4402] = 32'hFFFFFFF0;
    // rom_array[4403] = 32'hFFFFFFF0;
    // rom_array[4404] = 32'hFFFFFFF0;
    // rom_array[4405] = 32'h00002959;
    // rom_array[4406] = 32'hFFFFFFF0;
    // rom_array[4407] = 32'h00002961;
    // rom_array[4408] = 32'hFFFFFFF0;
    // rom_array[4409] = 32'hFFFFFFF0;
    // rom_array[4410] = 32'hFFFFFFF0;
    // rom_array[4411] = 32'hFFFFFFF0;
    // rom_array[4412] = 32'hFFFFFFF0;
    // rom_array[4413] = 32'h00002969;
    // rom_array[4414] = 32'hFFFFFFF0;
    // rom_array[4415] = 32'h00002971;
    // rom_array[4416] = 32'hFFFFFFF0;
    // rom_array[4417] = 32'hFFFFFFF1;
    // rom_array[4418] = 32'hFFFFFFF0;
    // rom_array[4419] = 32'hFFFFFFF1;
    // rom_array[4420] = 32'hFFFFFFF0;
    // rom_array[4421] = 32'h00002979;
    // rom_array[4422] = 32'hFFFFFFF0;
    // rom_array[4423] = 32'h00002981;
    // rom_array[4424] = 32'hFFFFFFF0;
    // rom_array[4425] = 32'hFFFFFFF1;
    // rom_array[4426] = 32'hFFFFFFF0;
    // rom_array[4427] = 32'hFFFFFFF1;
    // rom_array[4428] = 32'hFFFFFFF0;
    // rom_array[4429] = 32'h00002989;
    // rom_array[4430] = 32'hFFFFFFF0;
    // rom_array[4431] = 32'h00002991;
    // rom_array[4432] = 32'hFFFFFFF0;
    // rom_array[4433] = 32'hFFFFFFF0;
    // rom_array[4434] = 32'hFFFFFFF0;
    // rom_array[4435] = 32'hFFFFFFF0;
    // rom_array[4436] = 32'hFFFFFFF0;
    // rom_array[4437] = 32'h00002999;
    // rom_array[4438] = 32'hFFFFFFF0;
    // rom_array[4439] = 32'h000029a1;
    // rom_array[4440] = 32'hFFFFFFF0;
    // rom_array[4441] = 32'h000029a9;
    // rom_array[4442] = 32'hFFFFFFF0;
    // rom_array[4443] = 32'h000029b1;
    // rom_array[4444] = 32'hFFFFFFF0;
    // rom_array[4445] = 32'h000029b9;
    // rom_array[4446] = 32'hFFFFFFF0;
    // rom_array[4447] = 32'h000029c1;
    // rom_array[4448] = 32'hFFFFFFF0;
    // rom_array[4449] = 32'hFFFFFFF0;
    // rom_array[4450] = 32'hFFFFFFF0;
    // rom_array[4451] = 32'hFFFFFFF0;
    // rom_array[4452] = 32'hFFFFFFF0;
    // rom_array[4453] = 32'h000029c9;
    // rom_array[4454] = 32'hFFFFFFF0;
    // rom_array[4455] = 32'h000029d1;
    // rom_array[4456] = 32'hFFFFFFF0;
    // rom_array[4457] = 32'h000029d9;
    // rom_array[4458] = 32'hFFFFFFF0;
    // rom_array[4459] = 32'hFFFFFFF1;
    // rom_array[4460] = 32'hFFFFFFF0;
    // rom_array[4461] = 32'h000029e1;
    // rom_array[4462] = 32'hFFFFFFF0;
    // rom_array[4463] = 32'h000029e9;
    // rom_array[4464] = 32'hFFFFFFF0;
    // rom_array[4465] = 32'hFFFFFFF1;
    // rom_array[4466] = 32'hFFFFFFF0;
    // rom_array[4467] = 32'hFFFFFFF1;
    // rom_array[4468] = 32'hFFFFFFF0;
    // rom_array[4469] = 32'hFFFFFFF1;
    // rom_array[4470] = 32'hFFFFFFF0;
    // rom_array[4471] = 32'hFFFFFFF1;
    // rom_array[4472] = 32'hFFFFFFF0;
    // rom_array[4473] = 32'h000029f1;
    // rom_array[4474] = 32'hFFFFFFF0;
    // rom_array[4475] = 32'h000029f9;
    // rom_array[4476] = 32'hFFFFFFF0;
    // rom_array[4477] = 32'h00002a01;
    // rom_array[4478] = 32'hFFFFFFF0;
    // rom_array[4479] = 32'h00002a09;
    // rom_array[4480] = 32'hFFFFFFF0;
    // rom_array[4481] = 32'h00002a11;
    // rom_array[4482] = 32'hFFFFFFF0;
    // rom_array[4483] = 32'h00002a19;
    // rom_array[4484] = 32'hFFFFFFF0;
    // rom_array[4485] = 32'hFFFFFFF0;
    // rom_array[4486] = 32'hFFFFFFF0;
    // rom_array[4487] = 32'hFFFFFFF0;
    // rom_array[4488] = 32'hFFFFFFF0;
    // rom_array[4489] = 32'h00002a21;
    // rom_array[4490] = 32'hFFFFFFF0;
    // rom_array[4491] = 32'h00002a29;
    // rom_array[4492] = 32'hFFFFFFF0;
    // rom_array[4493] = 32'hFFFFFFF0;
    // rom_array[4494] = 32'hFFFFFFF0;
    // rom_array[4495] = 32'hFFFFFFF0;
    // rom_array[4496] = 32'hFFFFFFF0;
    // rom_array[4497] = 32'h00002a31;
    // rom_array[4498] = 32'hFFFFFFF0;
    // rom_array[4499] = 32'h00002a39;
    // rom_array[4500] = 32'hFFFFFFF0;
    // rom_array[4501] = 32'hFFFFFFF0;
    // rom_array[4502] = 32'hFFFFFFF0;
    // rom_array[4503] = 32'hFFFFFFF0;
    // rom_array[4504] = 32'hFFFFFFF0;
    // rom_array[4505] = 32'h00002a41;
    // rom_array[4506] = 32'hFFFFFFF0;
    // rom_array[4507] = 32'h00002a49;
    // rom_array[4508] = 32'hFFFFFFF0;
    // rom_array[4509] = 32'h00002a51;
    // rom_array[4510] = 32'hFFFFFFF0;
    // rom_array[4511] = 32'hFFFFFFF1;
    // rom_array[4512] = 32'hFFFFFFF0;
    // rom_array[4513] = 32'h00002a59;
    // rom_array[4514] = 32'hFFFFFFF0;
    // rom_array[4515] = 32'hFFFFFFF1;
    // rom_array[4516] = 32'hFFFFFFF0;
    // rom_array[4517] = 32'h00002a61;
    // rom_array[4518] = 32'hFFFFFFF0;
    // rom_array[4519] = 32'hFFFFFFF1;
    // rom_array[4520] = 32'hFFFFFFF0;
    // rom_array[4521] = 32'h00002a69;
    // rom_array[4522] = 32'hFFFFFFF0;
    // rom_array[4523] = 32'hFFFFFFF0;
    // rom_array[4524] = 32'hFFFFFFF0;
    // rom_array[4525] = 32'h00002a71;
    // rom_array[4526] = 32'hFFFFFFF0;
    // rom_array[4527] = 32'hFFFFFFF0;
    // rom_array[4528] = 32'hFFFFFFF0;
    // rom_array[4529] = 32'h00002a79;
    // rom_array[4530] = 32'hFFFFFFF0;
    // rom_array[4531] = 32'hFFFFFFF0;
    // rom_array[4532] = 32'hFFFFFFF0;
    // rom_array[4533] = 32'h00002a81;
    // rom_array[4534] = 32'hFFFFFFF0;
    // rom_array[4535] = 32'h00002a89;
    // rom_array[4536] = 32'hFFFFFFF0;
    // rom_array[4537] = 32'hFFFFFFF0;
    // rom_array[4538] = 32'hFFFFFFF0;
    // rom_array[4539] = 32'hFFFFFFF0;
    // rom_array[4540] = 32'hFFFFFFF0;
    // rom_array[4541] = 32'h00002a91;
    // rom_array[4542] = 32'hFFFFFFF0;
    // rom_array[4543] = 32'h00002a99;
    // rom_array[4544] = 32'hFFFFFFF0;
    // rom_array[4545] = 32'h00002aa1;
    // rom_array[4546] = 32'hFFFFFFF0;
    // rom_array[4547] = 32'hFFFFFFF1;
    // rom_array[4548] = 32'hFFFFFFF0;
    // rom_array[4549] = 32'h00002aa9;
    // rom_array[4550] = 32'hFFFFFFF0;
    // rom_array[4551] = 32'hFFFFFFF1;
    // rom_array[4552] = 32'hFFFFFFF0;
    // rom_array[4553] = 32'h00002ab1;
    // rom_array[4554] = 32'hFFFFFFF0;
    // rom_array[4555] = 32'hFFFFFFF1;
    // rom_array[4556] = 32'hFFFFFFF0;
    // rom_array[4557] = 32'h00002ab9;
    // rom_array[4558] = 32'hFFFFFFF0;
    // rom_array[4559] = 32'h00002ac1;
    // rom_array[4560] = 32'hFFFFFFF0;
    // rom_array[4561] = 32'h00002ac9;
    // rom_array[4562] = 32'hFFFFFFF0;
    // rom_array[4563] = 32'hFFFFFFF1;
    // rom_array[4564] = 32'hFFFFFFF0;
    // rom_array[4565] = 32'h00002ad1;
    // rom_array[4566] = 32'hFFFFFFF0;
    // rom_array[4567] = 32'h00002ad9;
    // rom_array[4568] = 32'hFFFFFFF0;
    // rom_array[4569] = 32'hFFFFFFF1;
    // rom_array[4570] = 32'hFFFFFFF0;
    // rom_array[4571] = 32'hFFFFFFF1;
    // rom_array[4572] = 32'hFFFFFFF0;
    // rom_array[4573] = 32'h00002ae1;
    // rom_array[4574] = 32'hFFFFFFF0;
    // rom_array[4575] = 32'h00002ae9;
    // rom_array[4576] = 32'hFFFFFFF0;
    // rom_array[4577] = 32'h00002af1;
    // rom_array[4578] = 32'hFFFFFFF0;
    // rom_array[4579] = 32'hFFFFFFF0;
    // rom_array[4580] = 32'hFFFFFFF0;
    // rom_array[4581] = 32'h00002af9;
    // rom_array[4582] = 32'hFFFFFFF0;
    // rom_array[4583] = 32'hFFFFFFF0;
    // rom_array[4584] = 32'hFFFFFFF0;
    // rom_array[4585] = 32'h00002b01;
    // rom_array[4586] = 32'hFFFFFFF0;
    // rom_array[4587] = 32'h00002b09;
    // rom_array[4588] = 32'hFFFFFFF0;
    // rom_array[4589] = 32'h00002b11;
    // rom_array[4590] = 32'hFFFFFFF0;
    // rom_array[4591] = 32'h00002b19;
    // rom_array[4592] = 32'hFFFFFFF0;
    // rom_array[4593] = 32'h00002b21;
    // rom_array[4594] = 32'hFFFFFFF0;
    // rom_array[4595] = 32'h00002b29;
    // rom_array[4596] = 32'hFFFFFFF0;
    // rom_array[4597] = 32'h00002b31;
    // rom_array[4598] = 32'hFFFFFFF0;
    // rom_array[4599] = 32'hFFFFFFF1;
    // rom_array[4600] = 32'hFFFFFFF0;
    // rom_array[4601] = 32'h00002b39;
    // rom_array[4602] = 32'hFFFFFFF0;
    // rom_array[4603] = 32'h00002b41;
    // rom_array[4604] = 32'hFFFFFFF0;
    // rom_array[4605] = 32'hFFFFFFF1;
    // rom_array[4606] = 32'hFFFFFFF0;
    // rom_array[4607] = 32'hFFFFFFF1;
    // rom_array[4608] = 32'hFFFFFFF0;
    // rom_array[4609] = 32'h00002b49;
    // rom_array[4610] = 32'hFFFFFFF0;
    // rom_array[4611] = 32'h00002b51;
    // rom_array[4612] = 32'hFFFFFFF0;
    // rom_array[4613] = 32'hFFFFFFF1;
    // rom_array[4614] = 32'hFFFFFFF0;
    // rom_array[4615] = 32'hFFFFFFF1;
    // rom_array[4616] = 32'hFFFFFFF0;
    // rom_array[4617] = 32'h00002b59;
    // rom_array[4618] = 32'hFFFFFFF0;
    // rom_array[4619] = 32'h00002b61;
    // rom_array[4620] = 32'hFFFFFFF0;
    // rom_array[4621] = 32'h00002b69;
    // rom_array[4622] = 32'hFFFFFFF0;
    // rom_array[4623] = 32'hFFFFFFF1;
    // rom_array[4624] = 32'hFFFFFFF0;
    // rom_array[4625] = 32'h00002b71;
    // rom_array[4626] = 32'hFFFFFFF0;
    // rom_array[4627] = 32'hFFFFFFF1;
    // rom_array[4628] = 32'hFFFFFFF0;
    // rom_array[4629] = 32'h00002b79;
    // rom_array[4630] = 32'hFFFFFFF0;
    // rom_array[4631] = 32'hFFFFFFF1;
    // rom_array[4632] = 32'hFFFFFFF0;
    // rom_array[4633] = 32'h00002b81;
    // rom_array[4634] = 32'hFFFFFFF0;
    // rom_array[4635] = 32'h00002b89;
    // rom_array[4636] = 32'hFFFFFFF0;
    // rom_array[4637] = 32'h00002b91;
    // rom_array[4638] = 32'hFFFFFFF0;
    // rom_array[4639] = 32'hFFFFFFF1;
    // rom_array[4640] = 32'hFFFFFFF0;
    // rom_array[4641] = 32'h00002b99;
    // rom_array[4642] = 32'hFFFFFFF0;
    // rom_array[4643] = 32'h00002ba1;
    // rom_array[4644] = 32'hFFFFFFF0;
    // rom_array[4645] = 32'h00002ba9;
    // rom_array[4646] = 32'hFFFFFFF0;
    // rom_array[4647] = 32'hFFFFFFF1;
    // rom_array[4648] = 32'hFFFFFFF0;
    // rom_array[4649] = 32'h00002bb1;
    // rom_array[4650] = 32'hFFFFFFF0;
    // rom_array[4651] = 32'h00002bb9;
    // rom_array[4652] = 32'hFFFFFFF0;
    // rom_array[4653] = 32'h00002bc1;
    // rom_array[4654] = 32'hFFFFFFF0;
    // rom_array[4655] = 32'hFFFFFFF1;
    // rom_array[4656] = 32'hFFFFFFF0;
    // rom_array[4657] = 32'h00002bc9;
    // rom_array[4658] = 32'hFFFFFFF0;
    // rom_array[4659] = 32'h00002bd1;
    // rom_array[4660] = 32'hFFFFFFF0;
    // rom_array[4661] = 32'h00002bd9;
    // rom_array[4662] = 32'hFFFFFFF0;
    // rom_array[4663] = 32'hFFFFFFF1;
    // rom_array[4664] = 32'hFFFFFFF0;
    // rom_array[4665] = 32'h00002be1;
    // rom_array[4666] = 32'hFFFFFFF0;
    // rom_array[4667] = 32'h00002be9;
    // rom_array[4668] = 32'hFFFFFFF0;
    // rom_array[4669] = 32'h00002bf1;
    // rom_array[4670] = 32'hFFFFFFF0;
    // rom_array[4671] = 32'h00002bf9;
    // rom_array[4672] = 32'hFFFFFFF0;
    // rom_array[4673] = 32'h00002c01;
    // rom_array[4674] = 32'hFFFFFFF0;
    // rom_array[4675] = 32'h00002c09;
    // rom_array[4676] = 32'hFFFFFFF0;
    // rom_array[4677] = 32'h00002c11;
    // rom_array[4678] = 32'hFFFFFFF0;
    // rom_array[4679] = 32'hFFFFFFF1;
    // rom_array[4680] = 32'hFFFFFFF0;
    // rom_array[4681] = 32'h00002c19;
    // rom_array[4682] = 32'hFFFFFFF0;
    // rom_array[4683] = 32'h00002c21;
    // rom_array[4684] = 32'hFFFFFFF0;
    // rom_array[4685] = 32'h00002c29;
    // rom_array[4686] = 32'hFFFFFFF0;
    // rom_array[4687] = 32'h00002c31;
    // rom_array[4688] = 32'hFFFFFFF0;
    // rom_array[4689] = 32'h00002c39;
    // rom_array[4690] = 32'hFFFFFFF0;
    // rom_array[4691] = 32'h00002c41;
    // rom_array[4692] = 32'hFFFFFFF0;
    // rom_array[4693] = 32'hFFFFFFF0;
    // rom_array[4694] = 32'hFFFFFFF0;
    // rom_array[4695] = 32'hFFFFFFF0;
    // rom_array[4696] = 32'hFFFFFFF0;
    // rom_array[4697] = 32'hFFFFFFF1;
    // rom_array[4698] = 32'hFFFFFFF0;
    // rom_array[4699] = 32'hFFFFFFF1;
    // rom_array[4700] = 32'hFFFFFFF0;
    // rom_array[4701] = 32'hFFFFFFF1;
    // rom_array[4702] = 32'hFFFFFFF0;
    // rom_array[4703] = 32'hFFFFFFF1;
    // rom_array[4704] = 32'hFFFFFFF0;
    // rom_array[4705] = 32'hFFFFFFF1;
    // rom_array[4706] = 32'hFFFFFFF0;
    // rom_array[4707] = 32'hFFFFFFF1;
    // rom_array[4708] = 32'hFFFFFFF0;
    // rom_array[4709] = 32'hFFFFFFF1;
    // rom_array[4710] = 32'hFFFFFFF0;
    // rom_array[4711] = 32'hFFFFFFF1;
    // rom_array[4712] = 32'hFFFFFFF0;
    // rom_array[4713] = 32'h00002c49;
    // rom_array[4714] = 32'hFFFFFFF0;
    // rom_array[4715] = 32'h00002c51;
    // rom_array[4716] = 32'hFFFFFFF0;
    // rom_array[4717] = 32'hFFFFFFF0;
    // rom_array[4718] = 32'hFFFFFFF0;
    // rom_array[4719] = 32'hFFFFFFF0;
    // rom_array[4720] = 32'hFFFFFFF0;
    // rom_array[4721] = 32'h00002c59;
    // rom_array[4722] = 32'hFFFFFFF0;
    // rom_array[4723] = 32'h00002c61;
    // rom_array[4724] = 32'hFFFFFFF0;
    // rom_array[4725] = 32'hFFFFFFF0;
    // rom_array[4726] = 32'hFFFFFFF0;
    // rom_array[4727] = 32'hFFFFFFF0;
    // rom_array[4728] = 32'hFFFFFFF0;
    // rom_array[4729] = 32'h00002c69;
    // rom_array[4730] = 32'hFFFFFFF0;
    // rom_array[4731] = 32'h00002c71;
    // rom_array[4732] = 32'hFFFFFFF0;
    // rom_array[4733] = 32'h00002c79;
    // rom_array[4734] = 32'hFFFFFFF0;
    // rom_array[4735] = 32'hFFFFFFF1;
    // rom_array[4736] = 32'hFFFFFFF0;
    // rom_array[4737] = 32'h00002c81;
    // rom_array[4738] = 32'hFFFFFFF0;
    // rom_array[4739] = 32'h00002c89;
    // rom_array[4740] = 32'hFFFFFFF0;
    // rom_array[4741] = 32'hFFFFFFF1;
    // rom_array[4742] = 32'hFFFFFFF0;
    // rom_array[4743] = 32'hFFFFFFF1;
    // rom_array[4744] = 32'hFFFFFFF0;
    // rom_array[4745] = 32'h00002c91;
    // rom_array[4746] = 32'hFFFFFFF0;
    // rom_array[4747] = 32'h00002c99;
    // rom_array[4748] = 32'hFFFFFFF0;
    // rom_array[4749] = 32'hFFFFFFF1;
    // rom_array[4750] = 32'hFFFFFFF0;
    // rom_array[4751] = 32'hFFFFFFF1;
    // rom_array[4752] = 32'hFFFFFFF0;
    // rom_array[4753] = 32'h00002ca1;
    // rom_array[4754] = 32'hFFFFFFF0;
    // rom_array[4755] = 32'h00002ca9;
    // rom_array[4756] = 32'hFFFFFFF0;
    // rom_array[4757] = 32'h00002cb1;
    // rom_array[4758] = 32'hFFFFFFF0;
    // rom_array[4759] = 32'hFFFFFFF1;
    // rom_array[4760] = 32'hFFFFFFF0;
    // rom_array[4761] = 32'h00002cb9;
    // rom_array[4762] = 32'hFFFFFFF0;
    // rom_array[4763] = 32'hFFFFFFF1;
    // rom_array[4764] = 32'hFFFFFFF0;
    // rom_array[4765] = 32'h00002cc1;
    // rom_array[4766] = 32'hFFFFFFF0;
    // rom_array[4767] = 32'hFFFFFFF1;
    // rom_array[4768] = 32'hFFFFFFF0;
    // rom_array[4769] = 32'h00002cc9;
    // rom_array[4770] = 32'hFFFFFFF0;
    // rom_array[4771] = 32'h00002cd1;
    // rom_array[4772] = 32'hFFFFFFF0;
    // rom_array[4773] = 32'h00002cd9;
    // rom_array[4774] = 32'hFFFFFFF0;
    // rom_array[4775] = 32'hFFFFFFF0;
    // rom_array[4776] = 32'hFFFFFFF0;
    // rom_array[4777] = 32'h00002ce1;
    // rom_array[4778] = 32'hFFFFFFF0;
    // rom_array[4779] = 32'h00002ce9;
    // rom_array[4780] = 32'hFFFFFFF0;
    // rom_array[4781] = 32'hFFFFFFF0;
    // rom_array[4782] = 32'hFFFFFFF0;
    // rom_array[4783] = 32'hFFFFFFF0;
    // rom_array[4784] = 32'hFFFFFFF0;
    // rom_array[4785] = 32'h00002cf1;
    // rom_array[4786] = 32'hFFFFFFF0;
    // rom_array[4787] = 32'hFFFFFFF0;
    // rom_array[4788] = 32'hFFFFFFF0;
    // rom_array[4789] = 32'h00002cf9;
    // rom_array[4790] = 32'hFFFFFFF0;
    // rom_array[4791] = 32'hFFFFFFF0;
    // rom_array[4792] = 32'hFFFFFFF0;
    // rom_array[4793] = 32'h00002d01;
    // rom_array[4794] = 32'hFFFFFFF0;
    // rom_array[4795] = 32'hFFFFFFF1;
    // rom_array[4796] = 32'hFFFFFFF0;
    // rom_array[4797] = 32'h00002d09;
    // rom_array[4798] = 32'hFFFFFFF0;
    // rom_array[4799] = 32'h00002d11;
    // rom_array[4800] = 32'hFFFFFFF0;
    // rom_array[4801] = 32'h00002d19;
    // rom_array[4802] = 32'hFFFFFFF0;
    // rom_array[4803] = 32'hFFFFFFF0;
    // rom_array[4804] = 32'hFFFFFFF0;
    // rom_array[4805] = 32'h00002d21;
    // rom_array[4806] = 32'hFFFFFFF0;
    // rom_array[4807] = 32'hFFFFFFF0;
    // rom_array[4808] = 32'hFFFFFFF0;
    // rom_array[4809] = 32'hFFFFFFF0;
    // rom_array[4810] = 32'h00002d29;
    // rom_array[4811] = 32'hFFFFFFF0;
    // rom_array[4812] = 32'hFFFFFFF0;
    // rom_array[4813] = 32'hFFFFFFF0;
    // rom_array[4814] = 32'hFFFFFFF0;
    // rom_array[4815] = 32'hFFFFFFF0;
    // rom_array[4816] = 32'hFFFFFFF0;
    // rom_array[4817] = 32'hFFFFFFF0;
    // rom_array[4818] = 32'hFFFFFFF0;
    // rom_array[4819] = 32'hFFFFFFF0;
    // rom_array[4820] = 32'h00002d31;
    // rom_array[4821] = 32'hFFFFFFF0;
    // rom_array[4822] = 32'hFFFFFFF0;
    // rom_array[4823] = 32'hFFFFFFF0;
    // rom_array[4824] = 32'hFFFFFFF0;
    // rom_array[4825] = 32'hFFFFFFF0;
    // rom_array[4826] = 32'h00002d39;
    // rom_array[4827] = 32'hFFFFFFF0;
    // rom_array[4828] = 32'h00002d41;
    // rom_array[4829] = 32'hFFFFFFF0;
    // rom_array[4830] = 32'hFFFFFFF0;
    // rom_array[4831] = 32'hFFFFFFF0;
    // rom_array[4832] = 32'hFFFFFFF0;
    // rom_array[4833] = 32'hFFFFFFF0;
    // rom_array[4834] = 32'hFFFFFFF0;
    // rom_array[4835] = 32'hFFFFFFF0;
    // rom_array[4836] = 32'hFFFFFFF0;
    // rom_array[4837] = 32'hFFFFFFF0;
    // rom_array[4838] = 32'h00002d49;
    // rom_array[4839] = 32'hFFFFFFF0;
    // rom_array[4840] = 32'h00002d51;
    // rom_array[4841] = 32'hFFFFFFF0;
    // rom_array[4842] = 32'hFFFFFFF0;
    // rom_array[4843] = 32'hFFFFFFF0;
    // rom_array[4844] = 32'hFFFFFFF0;
    // rom_array[4845] = 32'hFFFFFFF0;
    // rom_array[4846] = 32'h00002d59;
    // rom_array[4847] = 32'hFFFFFFF0;
    // rom_array[4848] = 32'h00002d61;
    // rom_array[4849] = 32'hFFFFFFF0;
    // rom_array[4850] = 32'hFFFFFFF1;
    // rom_array[4851] = 32'hFFFFFFF0;
    // rom_array[4852] = 32'hFFFFFFF1;
    // rom_array[4853] = 32'hFFFFFFF0;
    // rom_array[4854] = 32'h00002d69;
    // rom_array[4855] = 32'hFFFFFFF0;
    // rom_array[4856] = 32'h00002d71;
    // rom_array[4857] = 32'hFFFFFFF0;
    // rom_array[4858] = 32'hFFFFFFF1;
    // rom_array[4859] = 32'hFFFFFFF0;
    // rom_array[4860] = 32'hFFFFFFF1;
    // rom_array[4861] = 32'hFFFFFFF0;
    // rom_array[4862] = 32'h00002d79;
    // rom_array[4863] = 32'hFFFFFFF0;
    // rom_array[4864] = 32'h00002d81;
    // rom_array[4865] = 32'hFFFFFFF0;
    // rom_array[4866] = 32'hFFFFFFF0;
    // rom_array[4867] = 32'hFFFFFFF0;
    // rom_array[4868] = 32'hFFFFFFF0;
    // rom_array[4869] = 32'hFFFFFFF0;
    // rom_array[4870] = 32'h00002d89;
    // rom_array[4871] = 32'hFFFFFFF0;
    // rom_array[4872] = 32'h00002d91;
    // rom_array[4873] = 32'hFFFFFFF0;
    // rom_array[4874] = 32'hFFFFFFF1;
    // rom_array[4875] = 32'hFFFFFFF0;
    // rom_array[4876] = 32'h00002d99;
    // rom_array[4877] = 32'hFFFFFFF0;
    // rom_array[4878] = 32'h00002da1;
    // rom_array[4879] = 32'hFFFFFFF0;
    // rom_array[4880] = 32'h00002da9;
    // rom_array[4881] = 32'hFFFFFFF0;
    // rom_array[4882] = 32'h00002db1;
    // rom_array[4883] = 32'hFFFFFFF0;
    // rom_array[4884] = 32'hFFFFFFF0;
    // rom_array[4885] = 32'hFFFFFFF0;
    // rom_array[4886] = 32'h00002db9;
    // rom_array[4887] = 32'hFFFFFFF0;
    // rom_array[4888] = 32'hFFFFFFF0;
    // rom_array[4889] = 32'hFFFFFFF0;
    // rom_array[4890] = 32'hFFFFFFF0;
    // rom_array[4891] = 32'hFFFFFFF0;
    // rom_array[4892] = 32'h00002dc1;
    // rom_array[4893] = 32'hFFFFFFF0;
    // rom_array[4894] = 32'hFFFFFFF0;
    // rom_array[4895] = 32'hFFFFFFF0;
    // rom_array[4896] = 32'h00002dc9;
    // rom_array[4897] = 32'hFFFFFFF0;
    // rom_array[4898] = 32'h00002dd1;
    // rom_array[4899] = 32'hFFFFFFF0;
    // rom_array[4900] = 32'h00002dd9;
    // rom_array[4901] = 32'hFFFFFFF0;
    // rom_array[4902] = 32'h00002de1;
    // rom_array[4903] = 32'hFFFFFFF0;
    // rom_array[4904] = 32'hFFFFFFF1;
    // rom_array[4905] = 32'hFFFFFFF0;
    // rom_array[4906] = 32'h00002de9;
    // rom_array[4907] = 32'hFFFFFFF0;
    // rom_array[4908] = 32'h00002df1;
    // rom_array[4909] = 32'hFFFFFFF0;
    // rom_array[4910] = 32'hFFFFFFF1;
    // rom_array[4911] = 32'hFFFFFFF0;
    // rom_array[4912] = 32'h00002df9;
    // rom_array[4913] = 32'hFFFFFFF0;
    // rom_array[4914] = 32'hFFFFFFF1;
    // rom_array[4915] = 32'hFFFFFFF0;
    // rom_array[4916] = 32'h00002e01;
    // rom_array[4917] = 32'hFFFFFFF0;
    // rom_array[4918] = 32'hFFFFFFF1;
    // rom_array[4919] = 32'hFFFFFFF0;
    // rom_array[4920] = 32'h00002e09;
    // rom_array[4921] = 32'hFFFFFFF0;
    // rom_array[4922] = 32'hFFFFFFF1;
    // rom_array[4923] = 32'hFFFFFFF0;
    // rom_array[4924] = 32'h00002e11;
    // rom_array[4925] = 32'hFFFFFFF0;
    // rom_array[4926] = 32'h00002e19;
    // rom_array[4927] = 32'hFFFFFFF0;
    // rom_array[4928] = 32'h00002e21;
    // rom_array[4929] = 32'hFFFFFFF0;
    // rom_array[4930] = 32'h00002e29;
    // rom_array[4931] = 32'hFFFFFFF0;
    // rom_array[4932] = 32'h00002e31;
    // rom_array[4933] = 32'hFFFFFFF0;
    // rom_array[4934] = 32'hFFFFFFF0;
    // rom_array[4935] = 32'hFFFFFFF0;
    // rom_array[4936] = 32'hFFFFFFF0;
    // rom_array[4937] = 32'hFFFFFFF0;
    // rom_array[4938] = 32'h00002e39;
    // rom_array[4939] = 32'hFFFFFFF0;
    // rom_array[4940] = 32'h00002e41;
    // rom_array[4941] = 32'hFFFFFFF0;
    // rom_array[4942] = 32'hFFFFFFF0;
    // rom_array[4943] = 32'hFFFFFFF0;
    // rom_array[4944] = 32'hFFFFFFF0;
    // rom_array[4945] = 32'hFFFFFFF0;
    // rom_array[4946] = 32'hFFFFFFF0;
    // rom_array[4947] = 32'hFFFFFFF0;
    // rom_array[4948] = 32'h00002e49;
    // rom_array[4949] = 32'hFFFFFFF0;
    // rom_array[4950] = 32'hFFFFFFF0;
    // rom_array[4951] = 32'hFFFFFFF0;
    // rom_array[4952] = 32'h00002e51;
    // rom_array[4953] = 32'hFFFFFFF0;
    // rom_array[4954] = 32'hFFFFFFF0;
    // rom_array[4955] = 32'hFFFFFFF0;
    // rom_array[4956] = 32'hFFFFFFF0;
    // rom_array[4957] = 32'hFFFFFFF0;
    // rom_array[4958] = 32'h00002e59;
    // rom_array[4959] = 32'hFFFFFFF0;
    // rom_array[4960] = 32'h00002e61;
    // rom_array[4961] = 32'hFFFFFFF0;
    // rom_array[4962] = 32'hFFFFFFF0;
    // rom_array[4963] = 32'hFFFFFFF0;
    // rom_array[4964] = 32'h00002e69;
    // rom_array[4965] = 32'hFFFFFFF0;
    // rom_array[4966] = 32'h00002e71;
    // rom_array[4967] = 32'hFFFFFFF0;
    // rom_array[4968] = 32'h00002e79;
    // rom_array[4969] = 32'hFFFFFFF0;
    // rom_array[4970] = 32'h00002e81;
    // rom_array[4971] = 32'hFFFFFFF0;
    // rom_array[4972] = 32'h00002e89;
    // rom_array[4973] = 32'hFFFFFFF0;
    // rom_array[4974] = 32'hFFFFFFF1;
    // rom_array[4975] = 32'hFFFFFFF0;
    // rom_array[4976] = 32'h00002e91;
    // rom_array[4977] = 32'hFFFFFFF0;
    // rom_array[4978] = 32'hFFFFFFF1;
    // rom_array[4979] = 32'hFFFFFFF0;
    // rom_array[4980] = 32'h00002e99;
    // rom_array[4981] = 32'hFFFFFFF0;
    // rom_array[4982] = 32'hFFFFFFF1;
    // rom_array[4983] = 32'hFFFFFFF0;
    // rom_array[4984] = 32'h00002ea1;
    // rom_array[4985] = 32'hFFFFFFF0;
    // rom_array[4986] = 32'hFFFFFFF1;
    // rom_array[4987] = 32'hFFFFFFF0;
    // rom_array[4988] = 32'hFFFFFFF1;
    // rom_array[4989] = 32'hFFFFFFF0;
    // rom_array[4990] = 32'h00002ea9;
    // rom_array[4991] = 32'hFFFFFFF0;
    // rom_array[4992] = 32'h00002eb1;
    // rom_array[4993] = 32'hFFFFFFF0;
    // rom_array[4994] = 32'hFFFFFFF1;
    // rom_array[4995] = 32'hFFFFFFF0;
    // rom_array[4996] = 32'h00002eb9;
    // rom_array[4997] = 32'hFFFFFFF0;
    // rom_array[4998] = 32'h00002ec1;
    // rom_array[4999] = 32'hFFFFFFF0;
    // rom_array[5000] = 32'h00002ec9;
    // rom_array[5001] = 32'hFFFFFFF0;
    // rom_array[5002] = 32'hFFFFFFF0;
    // rom_array[5003] = 32'hFFFFFFF0;
    // rom_array[5004] = 32'h00002ed1;
    // rom_array[5005] = 32'hFFFFFFF0;
    // rom_array[5006] = 32'hFFFFFFF0;
    // rom_array[5007] = 32'hFFFFFFF0;
    // rom_array[5008] = 32'h00002ed9;
    // rom_array[5009] = 32'hFFFFFFF0;
    // rom_array[5010] = 32'hFFFFFFF1;
    // rom_array[5011] = 32'hFFFFFFF0;
    // rom_array[5012] = 32'h00002ee1;
    // rom_array[5013] = 32'hFFFFFFF0;
    // rom_array[5014] = 32'hFFFFFFF1;
    // rom_array[5015] = 32'hFFFFFFF0;
    // rom_array[5016] = 32'h00002ee9;
    // rom_array[5017] = 32'hFFFFFFF0;
    // rom_array[5018] = 32'hFFFFFFF1;
    // rom_array[5019] = 32'hFFFFFFF0;
    // rom_array[5020] = 32'h00002ef1;
    // rom_array[5021] = 32'hFFFFFFF0;
    // rom_array[5022] = 32'h00002ef9;
    // rom_array[5023] = 32'hFFFFFFF0;
    // rom_array[5024] = 32'h00002f01;
    // rom_array[5025] = 32'hFFFFFFF0;
    // rom_array[5026] = 32'h00002f09;
    // rom_array[5027] = 32'hFFFFFFF0;
    // rom_array[5028] = 32'h00002f11;
    // rom_array[5029] = 32'hFFFFFFF0;
    // rom_array[5030] = 32'hFFFFFFF1;
    // rom_array[5031] = 32'hFFFFFFF0;
    // rom_array[5032] = 32'hFFFFFFF1;
    // rom_array[5033] = 32'hFFFFFFF0;
    // rom_array[5034] = 32'h00002f19;
    // rom_array[5035] = 32'hFFFFFFF0;
    // rom_array[5036] = 32'h00002f21;
    // rom_array[5037] = 32'hFFFFFFF0;
    // rom_array[5038] = 32'hFFFFFFF1;
    // rom_array[5039] = 32'hFFFFFFF0;
    // rom_array[5040] = 32'hFFFFFFF1;
    // rom_array[5041] = 32'hFFFFFFF0;
    // rom_array[5042] = 32'hFFFFFFF1;
    // rom_array[5043] = 32'hFFFFFFF0;
    // rom_array[5044] = 32'hFFFFFFF1;
    // rom_array[5045] = 32'hFFFFFFF0;
    // rom_array[5046] = 32'hFFFFFFF1;
    // rom_array[5047] = 32'hFFFFFFF0;
    // rom_array[5048] = 32'hFFFFFFF1;
    // rom_array[5049] = 32'hFFFFFFF0;
    // rom_array[5050] = 32'hFFFFFFF1;
    // rom_array[5051] = 32'hFFFFFFF0;
    // rom_array[5052] = 32'hFFFFFFF1;
    // rom_array[5053] = 32'hFFFFFFF0;
    // rom_array[5054] = 32'hFFFFFFF1;
    // rom_array[5055] = 32'hFFFFFFF0;
    // rom_array[5056] = 32'hFFFFFFF1;
    // rom_array[5057] = 32'hFFFFFFF0;
    // rom_array[5058] = 32'h00002f29;
    // rom_array[5059] = 32'hFFFFFFF0;
    // rom_array[5060] = 32'h00002f31;
    // rom_array[5061] = 32'hFFFFFFF0;
    // rom_array[5062] = 32'hFFFFFFF1;
    // rom_array[5063] = 32'hFFFFFFF0;
    // rom_array[5064] = 32'h00002f39;
    // rom_array[5065] = 32'hFFFFFFF0;
    // rom_array[5066] = 32'hFFFFFFF1;
    // rom_array[5067] = 32'hFFFFFFF0;
    // rom_array[5068] = 32'h00002f41;
    // rom_array[5069] = 32'hFFFFFFF0;
    // rom_array[5070] = 32'hFFFFFFF1;
    // rom_array[5071] = 32'hFFFFFFF0;
    // rom_array[5072] = 32'h00002f49;
    // rom_array[5073] = 32'hFFFFFFF0;
    // rom_array[5074] = 32'h00002f51;
    // rom_array[5075] = 32'hFFFFFFF0;
    // rom_array[5076] = 32'h00002f59;
    // rom_array[5077] = 32'hFFFFFFF0;
    // rom_array[5078] = 32'hFFFFFFF1;
    // rom_array[5079] = 32'hFFFFFFF0;
    // rom_array[5080] = 32'hFFFFFFF1;
    // rom_array[5081] = 32'hFFFFFFF0;
    // rom_array[5082] = 32'h00002f61;
    // rom_array[5083] = 32'hFFFFFFF0;
    // rom_array[5084] = 32'h00002f69;
    // rom_array[5085] = 32'hFFFFFFF0;
    // rom_array[5086] = 32'hFFFFFFF1;
    // rom_array[5087] = 32'hFFFFFFF0;
    // rom_array[5088] = 32'h00002f71;
    // rom_array[5089] = 32'hFFFFFFF0;
    // rom_array[5090] = 32'h00002f79;
    // rom_array[5091] = 32'hFFFFFFF0;
    // rom_array[5092] = 32'h00002f81;
    // rom_array[5093] = 32'hFFFFFFF0;
    // rom_array[5094] = 32'hFFFFFFF1;
    // rom_array[5095] = 32'hFFFFFFF0;
    // rom_array[5096] = 32'hFFFFFFF1;
    // rom_array[5097] = 32'hFFFFFFF0;
    // rom_array[5098] = 32'h00002f89;
    // rom_array[5099] = 32'hFFFFFFF0;
    // rom_array[5100] = 32'h00002f91;
    // rom_array[5101] = 32'hFFFFFFF0;
    // rom_array[5102] = 32'hFFFFFFF1;
    // rom_array[5103] = 32'hFFFFFFF0;
    // rom_array[5104] = 32'hFFFFFFF1;
    // rom_array[5105] = 32'hFFFFFFF0;
    // rom_array[5106] = 32'h00002f99;
    // rom_array[5107] = 32'hFFFFFFF0;
    // rom_array[5108] = 32'h00002fa1;
    // rom_array[5109] = 32'hFFFFFFF0;
    // rom_array[5110] = 32'hFFFFFFF1;
    // rom_array[5111] = 32'hFFFFFFF0;
    // rom_array[5112] = 32'h00002fa9;
    // rom_array[5113] = 32'hFFFFFFF0;
    // rom_array[5114] = 32'h00002fb1;
    // rom_array[5115] = 32'hFFFFFFF0;
    // rom_array[5116] = 32'h00002fb9;
    // rom_array[5117] = 32'hFFFFFFF0;
    // rom_array[5118] = 32'hFFFFFFF1;
    // rom_array[5119] = 32'hFFFFFFF0;
    // rom_array[5120] = 32'h00002fc1;
    // rom_array[5121] = 32'hFFFFFFF0;
    // rom_array[5122] = 32'hFFFFFFF1;
    // rom_array[5123] = 32'hFFFFFFF0;
    // rom_array[5124] = 32'hFFFFFFF1;
    // rom_array[5125] = 32'hFFFFFFF0;
    // rom_array[5126] = 32'hFFFFFFF1;
    // rom_array[5127] = 32'hFFFFFFF0;
    // rom_array[5128] = 32'hFFFFFFF1;
    // rom_array[5129] = 32'hFFFFFFF0;
    // rom_array[5130] = 32'hFFFFFFF1;
    // rom_array[5131] = 32'hFFFFFFF0;
    // rom_array[5132] = 32'hFFFFFFF1;
    // rom_array[5133] = 32'hFFFFFFF0;
    // rom_array[5134] = 32'hFFFFFFF1;
    // rom_array[5135] = 32'hFFFFFFF0;
    // rom_array[5136] = 32'hFFFFFFF1;
    // rom_array[5137] = 32'hFFFFFFF0;
    // rom_array[5138] = 32'h00002fc9;
    // rom_array[5139] = 32'hFFFFFFF0;
    // rom_array[5140] = 32'h00002fd1;
    // rom_array[5141] = 32'hFFFFFFF0;
    // rom_array[5142] = 32'hFFFFFFF0;
    // rom_array[5143] = 32'hFFFFFFF0;
    // rom_array[5144] = 32'hFFFFFFF0;
    // rom_array[5145] = 32'hFFFFFFF0;
    // rom_array[5146] = 32'h00002fd9;
    // rom_array[5147] = 32'hFFFFFFF0;
    // rom_array[5148] = 32'h00002fe1;
    // rom_array[5149] = 32'hFFFFFFF0;
    // rom_array[5150] = 32'hFFFFFFF0;
    // rom_array[5151] = 32'hFFFFFFF0;
    // rom_array[5152] = 32'hFFFFFFF0;
    // rom_array[5153] = 32'hFFFFFFF0;
    // rom_array[5154] = 32'hFFFFFFF1;
    // rom_array[5155] = 32'hFFFFFFF0;
    // rom_array[5156] = 32'h00002fe9;
    // rom_array[5157] = 32'hFFFFFFF0;
    // rom_array[5158] = 32'hFFFFFFF1;
    // rom_array[5159] = 32'hFFFFFFF0;
    // rom_array[5160] = 32'h00002ff1;
    // rom_array[5161] = 32'hFFFFFFF0;
    // rom_array[5162] = 32'h00002ff9;
    // rom_array[5163] = 32'hFFFFFFF0;
    // rom_array[5164] = 32'h00003001;
    // rom_array[5165] = 32'hFFFFFFF0;
    // rom_array[5166] = 32'hFFFFFFF0;
    // rom_array[5167] = 32'hFFFFFFF0;
    // rom_array[5168] = 32'hFFFFFFF0;
    // rom_array[5169] = 32'hFFFFFFF0;
    // rom_array[5170] = 32'h00003009;
    // rom_array[5171] = 32'hFFFFFFF0;
    // rom_array[5172] = 32'h00003011;
    // rom_array[5173] = 32'hFFFFFFF0;
    // rom_array[5174] = 32'hFFFFFFF1;
    // rom_array[5175] = 32'hFFFFFFF0;
    // rom_array[5176] = 32'hFFFFFFF1;
    // rom_array[5177] = 32'hFFFFFFF0;
    // rom_array[5178] = 32'h00003019;
    // rom_array[5179] = 32'hFFFFFFF0;
    // rom_array[5180] = 32'h00003021;
    // rom_array[5181] = 32'hFFFFFFF0;
    // rom_array[5182] = 32'hFFFFFFF1;
    // rom_array[5183] = 32'hFFFFFFF0;
    // rom_array[5184] = 32'hFFFFFFF1;
    // rom_array[5185] = 32'hFFFFFFF0;
    // rom_array[5186] = 32'h00003029;
    // rom_array[5187] = 32'hFFFFFFF0;
    // rom_array[5188] = 32'h00003031;
    // rom_array[5189] = 32'hFFFFFFF0;
    // rom_array[5190] = 32'hFFFFFFF1;
    // rom_array[5191] = 32'hFFFFFFF0;
    // rom_array[5192] = 32'h00003039;
    // rom_array[5193] = 32'hFFFFFFF0;
    // rom_array[5194] = 32'h00003041;
    // rom_array[5195] = 32'hFFFFFFF0;
    // rom_array[5196] = 32'h00003049;
    // rom_array[5197] = 32'hFFFFFFF0;
    // rom_array[5198] = 32'hFFFFFFF0;
    // rom_array[5199] = 32'hFFFFFFF0;
    // rom_array[5200] = 32'hFFFFFFF0;
    // rom_array[5201] = 32'hFFFFFFF0;
    // rom_array[5202] = 32'h00003051;
    // rom_array[5203] = 32'hFFFFFFF0;
    // rom_array[5204] = 32'h00003059;
    // rom_array[5205] = 32'hFFFFFFF0;
    // rom_array[5206] = 32'hFFFFFFF0;
    // rom_array[5207] = 32'hFFFFFFF0;
    // rom_array[5208] = 32'hFFFFFFF0;
    // rom_array[5209] = 32'hFFFFFFF0;
    // rom_array[5210] = 32'h00003061;
    // rom_array[5211] = 32'hFFFFFFF0;
    // rom_array[5212] = 32'h00003069;
    // rom_array[5213] = 32'hFFFFFFF0;
    // rom_array[5214] = 32'hFFFFFFF0;
    // rom_array[5215] = 32'hFFFFFFF0;
    // rom_array[5216] = 32'hFFFFFFF0;
    // rom_array[5217] = 32'h00003071;
    // rom_array[5218] = 32'hFFFFFFF0;
    // rom_array[5219] = 32'hFFFFFFF0;
    // rom_array[5220] = 32'hFFFFFFF0;
    // rom_array[5221] = 32'hFFFFFFF0;
    // rom_array[5222] = 32'hFFFFFFF0;
    // rom_array[5223] = 32'hFFFFFFF0;
    // rom_array[5224] = 32'hFFFFFFF0;
    // rom_array[5225] = 32'hFFFFFFF0;
    // rom_array[5226] = 32'hFFFFFFF0;
    // rom_array[5227] = 32'h00003079;
    // rom_array[5228] = 32'hFFFFFFF0;
    // rom_array[5229] = 32'hFFFFFFF0;
    // rom_array[5230] = 32'hFFFFFFF0;
    // rom_array[5231] = 32'hFFFFFFF0;
    // rom_array[5232] = 32'hFFFFFFF0;
    // rom_array[5233] = 32'h00003081;
    // rom_array[5234] = 32'hFFFFFFF0;
    // rom_array[5235] = 32'h00003089;
    // rom_array[5236] = 32'hFFFFFFF0;
    // rom_array[5237] = 32'hFFFFFFF0;
    // rom_array[5238] = 32'hFFFFFFF0;
    // rom_array[5239] = 32'hFFFFFFF0;
    // rom_array[5240] = 32'hFFFFFFF0;
    // rom_array[5241] = 32'hFFFFFFF0;
    // rom_array[5242] = 32'hFFFFFFF0;
    // rom_array[5243] = 32'hFFFFFFF0;
    // rom_array[5244] = 32'hFFFFFFF0;
    // rom_array[5245] = 32'h00003091;
    // rom_array[5246] = 32'hFFFFFFF0;
    // rom_array[5247] = 32'h00003099;
    // rom_array[5248] = 32'hFFFFFFF0;
    // rom_array[5249] = 32'hFFFFFFF0;
    // rom_array[5250] = 32'hFFFFFFF0;
    // rom_array[5251] = 32'hFFFFFFF0;
    // rom_array[5252] = 32'hFFFFFFF0;
    // rom_array[5253] = 32'h000030a1;
    // rom_array[5254] = 32'hFFFFFFF0;
    // rom_array[5255] = 32'h000030a9;
    // rom_array[5256] = 32'hFFFFFFF0;
    // rom_array[5257] = 32'hFFFFFFF1;
    // rom_array[5258] = 32'hFFFFFFF0;
    // rom_array[5259] = 32'hFFFFFFF1;
    // rom_array[5260] = 32'hFFFFFFF0;
    // rom_array[5261] = 32'h000030b1;
    // rom_array[5262] = 32'hFFFFFFF0;
    // rom_array[5263] = 32'h000030b9;
    // rom_array[5264] = 32'hFFFFFFF0;
    // rom_array[5265] = 32'hFFFFFFF1;
    // rom_array[5266] = 32'hFFFFFFF0;
    // rom_array[5267] = 32'hFFFFFFF1;
    // rom_array[5268] = 32'hFFFFFFF0;
    // rom_array[5269] = 32'h000030c1;
    // rom_array[5270] = 32'hFFFFFFF0;
    // rom_array[5271] = 32'h000030c9;
    // rom_array[5272] = 32'hFFFFFFF0;
    // rom_array[5273] = 32'hFFFFFFF0;
    // rom_array[5274] = 32'hFFFFFFF0;
    // rom_array[5275] = 32'hFFFFFFF0;
    // rom_array[5276] = 32'hFFFFFFF0;
    // rom_array[5277] = 32'h000030d1;
    // rom_array[5278] = 32'hFFFFFFF0;
    // rom_array[5279] = 32'h000030d9;
    // rom_array[5280] = 32'hFFFFFFF0;
    // rom_array[5281] = 32'hFFFFFFF1;
    // rom_array[5282] = 32'hFFFFFFF0;
    // rom_array[5283] = 32'h000030e1;
    // rom_array[5284] = 32'hFFFFFFF0;
    // rom_array[5285] = 32'h000030e9;
    // rom_array[5286] = 32'hFFFFFFF0;
    // rom_array[5287] = 32'h000030f1;
    // rom_array[5288] = 32'hFFFFFFF0;
    // rom_array[5289] = 32'h000030f9;
    // rom_array[5290] = 32'hFFFFFFF0;
    // rom_array[5291] = 32'hFFFFFFF0;
    // rom_array[5292] = 32'hFFFFFFF0;
    // rom_array[5293] = 32'h00003101;
    // rom_array[5294] = 32'hFFFFFFF0;
    // rom_array[5295] = 32'hFFFFFFF0;
    // rom_array[5296] = 32'hFFFFFFF0;
    // rom_array[5297] = 32'hFFFFFFF0;
    // rom_array[5298] = 32'hFFFFFFF0;
    // rom_array[5299] = 32'h00003109;
    // rom_array[5300] = 32'hFFFFFFF0;
    // rom_array[5301] = 32'hFFFFFFF0;
    // rom_array[5302] = 32'hFFFFFFF0;
    // rom_array[5303] = 32'h00003111;
    // rom_array[5304] = 32'hFFFFFFF0;
    // rom_array[5305] = 32'h00003119;
    // rom_array[5306] = 32'hFFFFFFF0;
    // rom_array[5307] = 32'h00003121;
    // rom_array[5308] = 32'hFFFFFFF0;
    // rom_array[5309] = 32'h00003129;
    // rom_array[5310] = 32'hFFFFFFF0;
    // rom_array[5311] = 32'hFFFFFFF1;
    // rom_array[5312] = 32'hFFFFFFF0;
    // rom_array[5313] = 32'h00003131;
    // rom_array[5314] = 32'hFFFFFFF0;
    // rom_array[5315] = 32'h00003139;
    // rom_array[5316] = 32'hFFFFFFF0;
    // rom_array[5317] = 32'hFFFFFFF1;
    // rom_array[5318] = 32'hFFFFFFF0;
    // rom_array[5319] = 32'h00003141;
    // rom_array[5320] = 32'hFFFFFFF0;
    // rom_array[5321] = 32'hFFFFFFF1;
    // rom_array[5322] = 32'hFFFFFFF0;
    // rom_array[5323] = 32'h00003149;
    // rom_array[5324] = 32'hFFFFFFF0;
    // rom_array[5325] = 32'hFFFFFFF1;
    // rom_array[5326] = 32'hFFFFFFF0;
    // rom_array[5327] = 32'h00003151;
    // rom_array[5328] = 32'hFFFFFFF0;
    // rom_array[5329] = 32'hFFFFFFF1;
    // rom_array[5330] = 32'hFFFFFFF0;
    // rom_array[5331] = 32'h00003159;
    // rom_array[5332] = 32'hFFFFFFF0;
    // rom_array[5333] = 32'h00003161;
    // rom_array[5334] = 32'hFFFFFFF0;
    // rom_array[5335] = 32'h00003169;
    // rom_array[5336] = 32'hFFFFFFF0;
    // rom_array[5337] = 32'h00003171;
    // rom_array[5338] = 32'hFFFFFFF0;
    // rom_array[5339] = 32'h00003179;
    // rom_array[5340] = 32'hFFFFFFF0;
    // rom_array[5341] = 32'hFFFFFFF0;
    // rom_array[5342] = 32'hFFFFFFF0;
    // rom_array[5343] = 32'hFFFFFFF0;
    // rom_array[5344] = 32'hFFFFFFF0;
    // rom_array[5345] = 32'h00003181;
    // rom_array[5346] = 32'hFFFFFFF0;
    // rom_array[5347] = 32'h00003189;
    // rom_array[5348] = 32'hFFFFFFF0;
    // rom_array[5349] = 32'hFFFFFFF0;
    // rom_array[5350] = 32'hFFFFFFF0;
    // rom_array[5351] = 32'hFFFFFFF0;
    // rom_array[5352] = 32'hFFFFFFF0;
    // rom_array[5353] = 32'hFFFFFFF0;
    // rom_array[5354] = 32'hFFFFFFF0;
    // rom_array[5355] = 32'h00003191;
    // rom_array[5356] = 32'hFFFFFFF0;
    // rom_array[5357] = 32'hFFFFFFF0;
    // rom_array[5358] = 32'hFFFFFFF0;
    // rom_array[5359] = 32'h00003199;
    // rom_array[5360] = 32'hFFFFFFF0;
    // rom_array[5361] = 32'hFFFFFFF0;
    // rom_array[5362] = 32'hFFFFFFF0;
    // rom_array[5363] = 32'hFFFFFFF0;
    // rom_array[5364] = 32'hFFFFFFF0;
    // rom_array[5365] = 32'h000031a1;
    // rom_array[5366] = 32'hFFFFFFF0;
    // rom_array[5367] = 32'h000031a9;
    // rom_array[5368] = 32'hFFFFFFF0;
    // rom_array[5369] = 32'hFFFFFFF0;
    // rom_array[5370] = 32'hFFFFFFF0;
    // rom_array[5371] = 32'h000031b1;
    // rom_array[5372] = 32'hFFFFFFF0;
    // rom_array[5373] = 32'h000031b9;
    // rom_array[5374] = 32'hFFFFFFF0;
    // rom_array[5375] = 32'h000031c1;
    // rom_array[5376] = 32'hFFFFFFF0;
    // rom_array[5377] = 32'h000031c9;
    // rom_array[5378] = 32'hFFFFFFF0;
    // rom_array[5379] = 32'h000031d1;
    // rom_array[5380] = 32'hFFFFFFF0;
    // rom_array[5381] = 32'hFFFFFFF1;
    // rom_array[5382] = 32'hFFFFFFF0;
    // rom_array[5383] = 32'h000031d9;
    // rom_array[5384] = 32'hFFFFFFF0;
    // rom_array[5385] = 32'hFFFFFFF1;
    // rom_array[5386] = 32'hFFFFFFF0;
    // rom_array[5387] = 32'h000031e1;
    // rom_array[5388] = 32'hFFFFFFF0;
    // rom_array[5389] = 32'hFFFFFFF1;
    // rom_array[5390] = 32'hFFFFFFF0;
    // rom_array[5391] = 32'h000031e9;
    // rom_array[5392] = 32'hFFFFFFF0;
    // rom_array[5393] = 32'hFFFFFFF1;
    // rom_array[5394] = 32'hFFFFFFF0;
    // rom_array[5395] = 32'hFFFFFFF1;
    // rom_array[5396] = 32'hFFFFFFF0;
    // rom_array[5397] = 32'h000031f1;
    // rom_array[5398] = 32'hFFFFFFF0;
    // rom_array[5399] = 32'h000031f9;
    // rom_array[5400] = 32'hFFFFFFF0;
    // rom_array[5401] = 32'hFFFFFFF1;
    // rom_array[5402] = 32'hFFFFFFF0;
    // rom_array[5403] = 32'h00003201;
    // rom_array[5404] = 32'hFFFFFFF0;
    // rom_array[5405] = 32'h00003209;
    // rom_array[5406] = 32'hFFFFFFF0;
    // rom_array[5407] = 32'h00003211;
    // rom_array[5408] = 32'hFFFFFFF0;
    // rom_array[5409] = 32'hFFFFFFF0;
    // rom_array[5410] = 32'hFFFFFFF0;
    // rom_array[5411] = 32'h00003219;
    // rom_array[5412] = 32'hFFFFFFF0;
    // rom_array[5413] = 32'hFFFFFFF0;
    // rom_array[5414] = 32'hFFFFFFF0;
    // rom_array[5415] = 32'h00003221;
    // rom_array[5416] = 32'hFFFFFFF0;
    // rom_array[5417] = 32'hFFFFFFF1;
    // rom_array[5418] = 32'hFFFFFFF0;
    // rom_array[5419] = 32'h00003229;
    // rom_array[5420] = 32'hFFFFFFF0;
    // rom_array[5421] = 32'hFFFFFFF1;
    // rom_array[5422] = 32'hFFFFFFF0;
    // rom_array[5423] = 32'h00003231;
    // rom_array[5424] = 32'hFFFFFFF0;
    // rom_array[5425] = 32'hFFFFFFF1;
    // rom_array[5426] = 32'hFFFFFFF0;
    // rom_array[5427] = 32'h00003239;
    // rom_array[5428] = 32'hFFFFFFF0;
    // rom_array[5429] = 32'h00003241;
    // rom_array[5430] = 32'hFFFFFFF0;
    // rom_array[5431] = 32'h00003249;
    // rom_array[5432] = 32'hFFFFFFF0;
    // rom_array[5433] = 32'h00003251;
    // rom_array[5434] = 32'hFFFFFFF0;
    // rom_array[5435] = 32'h00003259;
    // rom_array[5436] = 32'hFFFFFFF0;
    // rom_array[5437] = 32'hFFFFFFF1;
    // rom_array[5438] = 32'hFFFFFFF0;
    // rom_array[5439] = 32'hFFFFFFF1;
    // rom_array[5440] = 32'hFFFFFFF0;
    // rom_array[5441] = 32'h00003261;
    // rom_array[5442] = 32'hFFFFFFF0;
    // rom_array[5443] = 32'h00003269;
    // rom_array[5444] = 32'hFFFFFFF0;
    // rom_array[5445] = 32'hFFFFFFF1;
    // rom_array[5446] = 32'hFFFFFFF0;
    // rom_array[5447] = 32'hFFFFFFF1;
    // rom_array[5448] = 32'hFFFFFFF0;
    // rom_array[5449] = 32'hFFFFFFF1;
    // rom_array[5450] = 32'hFFFFFFF0;
    // rom_array[5451] = 32'hFFFFFFF1;
    // rom_array[5452] = 32'hFFFFFFF0;
    // rom_array[5453] = 32'hFFFFFFF1;
    // rom_array[5454] = 32'hFFFFFFF0;
    // rom_array[5455] = 32'hFFFFFFF1;
    // rom_array[5456] = 32'hFFFFFFF0;
    // rom_array[5457] = 32'hFFFFFFF1;
    // rom_array[5458] = 32'hFFFFFFF0;
    // rom_array[5459] = 32'hFFFFFFF1;
    // rom_array[5460] = 32'hFFFFFFF0;
    // rom_array[5461] = 32'hFFFFFFF1;
    // rom_array[5462] = 32'hFFFFFFF0;
    // rom_array[5463] = 32'hFFFFFFF1;
    // rom_array[5464] = 32'hFFFFFFF0;
    // rom_array[5465] = 32'h00003271;
    // rom_array[5466] = 32'hFFFFFFF0;
    // rom_array[5467] = 32'h00003279;
    // rom_array[5468] = 32'hFFFFFFF0;
    // rom_array[5469] = 32'hFFFFFFF1;
    // rom_array[5470] = 32'hFFFFFFF0;
    // rom_array[5471] = 32'h00003281;
    // rom_array[5472] = 32'hFFFFFFF0;
    // rom_array[5473] = 32'hFFFFFFF1;
    // rom_array[5474] = 32'hFFFFFFF0;
    // rom_array[5475] = 32'h00003289;
    // rom_array[5476] = 32'hFFFFFFF0;
    // rom_array[5477] = 32'hFFFFFFF1;
    // rom_array[5478] = 32'hFFFFFFF0;
    // rom_array[5479] = 32'h00003291;
    // rom_array[5480] = 32'hFFFFFFF0;
    // rom_array[5481] = 32'h00003299;
    // rom_array[5482] = 32'hFFFFFFF0;
    // rom_array[5483] = 32'h000032a1;
    // rom_array[5484] = 32'hFFFFFFF0;
    // rom_array[5485] = 32'hFFFFFFF1;
    // rom_array[5486] = 32'hFFFFFFF0;
    // rom_array[5487] = 32'hFFFFFFF1;
    // rom_array[5488] = 32'hFFFFFFF0;
    // rom_array[5489] = 32'h000032a9;
    // rom_array[5490] = 32'hFFFFFFF0;
    // rom_array[5491] = 32'h000032b1;
    // rom_array[5492] = 32'hFFFFFFF0;
    // rom_array[5493] = 32'hFFFFFFF1;
    // rom_array[5494] = 32'hFFFFFFF0;
    // rom_array[5495] = 32'h000032b9;
    // rom_array[5496] = 32'hFFFFFFF0;
    // rom_array[5497] = 32'h000032c1;
    // rom_array[5498] = 32'hFFFFFFF0;
    // rom_array[5499] = 32'h000032c9;
    // rom_array[5500] = 32'hFFFFFFF0;
    // rom_array[5501] = 32'hFFFFFFF1;
    // rom_array[5502] = 32'hFFFFFFF0;
    // rom_array[5503] = 32'hFFFFFFF1;
    // rom_array[5504] = 32'hFFFFFFF0;
    // rom_array[5505] = 32'h000032d1;
    // rom_array[5506] = 32'hFFFFFFF0;
    // rom_array[5507] = 32'h000032d9;
    // rom_array[5508] = 32'hFFFFFFF0;
    // rom_array[5509] = 32'hFFFFFFF1;
    // rom_array[5510] = 32'hFFFFFFF0;
    // rom_array[5511] = 32'hFFFFFFF1;
    // rom_array[5512] = 32'hFFFFFFF0;
    // rom_array[5513] = 32'h000032e1;
    // rom_array[5514] = 32'hFFFFFFF0;
    // rom_array[5515] = 32'h000032e9;
    // rom_array[5516] = 32'hFFFFFFF0;
    // rom_array[5517] = 32'hFFFFFFF1;
    // rom_array[5518] = 32'hFFFFFFF0;
    // rom_array[5519] = 32'h000032f1;
    // rom_array[5520] = 32'hFFFFFFF0;
    // rom_array[5521] = 32'h000032f9;
    // rom_array[5522] = 32'hFFFFFFF0;
    // rom_array[5523] = 32'h00003301;
    // rom_array[5524] = 32'hFFFFFFF0;
    // rom_array[5525] = 32'hFFFFFFF1;
    // rom_array[5526] = 32'hFFFFFFF0;
    // rom_array[5527] = 32'h00003309;
    // rom_array[5528] = 32'hFFFFFFF0;
    // rom_array[5529] = 32'hFFFFFFF1;
    // rom_array[5530] = 32'hFFFFFFF0;
    // rom_array[5531] = 32'hFFFFFFF1;
    // rom_array[5532] = 32'hFFFFFFF0;
    // rom_array[5533] = 32'hFFFFFFF1;
    // rom_array[5534] = 32'hFFFFFFF0;
    // rom_array[5535] = 32'hFFFFFFF1;
    // rom_array[5536] = 32'hFFFFFFF0;
    // rom_array[5537] = 32'hFFFFFFF1;
    // rom_array[5538] = 32'hFFFFFFF0;
    // rom_array[5539] = 32'hFFFFFFF1;
    // rom_array[5540] = 32'hFFFFFFF0;
    // rom_array[5541] = 32'hFFFFFFF1;
    // rom_array[5542] = 32'hFFFFFFF0;
    // rom_array[5543] = 32'hFFFFFFF1;
    // rom_array[5544] = 32'hFFFFFFF0;
    // rom_array[5545] = 32'h00003311;
    // rom_array[5546] = 32'hFFFFFFF0;
    // rom_array[5547] = 32'h00003319;
    // rom_array[5548] = 32'hFFFFFFF0;
    // rom_array[5549] = 32'hFFFFFFF0;
    // rom_array[5550] = 32'hFFFFFFF0;
    // rom_array[5551] = 32'hFFFFFFF0;
    // rom_array[5552] = 32'hFFFFFFF0;
    // rom_array[5553] = 32'h00003321;
    // rom_array[5554] = 32'hFFFFFFF0;
    // rom_array[5555] = 32'h00003329;
    // rom_array[5556] = 32'hFFFFFFF0;
    // rom_array[5557] = 32'hFFFFFFF0;
    // rom_array[5558] = 32'hFFFFFFF0;
    // rom_array[5559] = 32'hFFFFFFF0;
    // rom_array[5560] = 32'hFFFFFFF0;
    // rom_array[5561] = 32'hFFFFFFF1;
    // rom_array[5562] = 32'hFFFFFFF0;
    // rom_array[5563] = 32'h00003331;
    // rom_array[5564] = 32'hFFFFFFF0;
    // rom_array[5565] = 32'hFFFFFFF1;
    // rom_array[5566] = 32'hFFFFFFF0;
    // rom_array[5567] = 32'h00003339;
    // rom_array[5568] = 32'hFFFFFFF0;
    // rom_array[5569] = 32'h00003341;
    // rom_array[5570] = 32'hFFFFFFF0;
    // rom_array[5571] = 32'h00003349;
    // rom_array[5572] = 32'hFFFFFFF0;
    // rom_array[5573] = 32'hFFFFFFF0;
    // rom_array[5574] = 32'hFFFFFFF0;
    // rom_array[5575] = 32'hFFFFFFF0;
    // rom_array[5576] = 32'hFFFFFFF0;
    // rom_array[5577] = 32'h00003351;
    // rom_array[5578] = 32'hFFFFFFF0;
    // rom_array[5579] = 32'h00003359;
    // rom_array[5580] = 32'hFFFFFFF0;
    // rom_array[5581] = 32'hFFFFFFF1;
    // rom_array[5582] = 32'hFFFFFFF0;
    // rom_array[5583] = 32'hFFFFFFF1;
    // rom_array[5584] = 32'hFFFFFFF0;
    // rom_array[5585] = 32'h00003361;
    // rom_array[5586] = 32'hFFFFFFF0;
    // rom_array[5587] = 32'h00003369;
    // rom_array[5588] = 32'hFFFFFFF0;
    // rom_array[5589] = 32'hFFFFFFF1;
    // rom_array[5590] = 32'hFFFFFFF0;
    // rom_array[5591] = 32'hFFFFFFF1;
    // rom_array[5592] = 32'hFFFFFFF0;
    // rom_array[5593] = 32'h00003371;
    // rom_array[5594] = 32'hFFFFFFF0;
    // rom_array[5595] = 32'h00003379;
    // rom_array[5596] = 32'hFFFFFFF0;
    // rom_array[5597] = 32'hFFFFFFF1;
    // rom_array[5598] = 32'hFFFFFFF0;
    // rom_array[5599] = 32'h00003381;
    // rom_array[5600] = 32'hFFFFFFF0;
    // rom_array[5601] = 32'h00003389;
    // rom_array[5602] = 32'hFFFFFFF0;
    // rom_array[5603] = 32'h00003391;
    // rom_array[5604] = 32'hFFFFFFF0;
    // rom_array[5605] = 32'hFFFFFFF0;
    // rom_array[5606] = 32'hFFFFFFF0;
    // rom_array[5607] = 32'hFFFFFFF0;
    // rom_array[5608] = 32'hFFFFFFF0;
    // rom_array[5609] = 32'h00003399;
    // rom_array[5610] = 32'hFFFFFFF0;
    // rom_array[5611] = 32'h000033a1;
    // rom_array[5612] = 32'hFFFFFFF0;
    // rom_array[5613] = 32'hFFFFFFF0;
    // rom_array[5614] = 32'hFFFFFFF0;
    // rom_array[5615] = 32'hFFFFFFF0;
    // rom_array[5616] = 32'hFFFFFFF0;
    // rom_array[5617] = 32'h000033a9;
    // rom_array[5618] = 32'hFFFFFFF0;
    // rom_array[5619] = 32'h000033b1;
    // rom_array[5620] = 32'hFFFFFFF0;
    // rom_array[5621] = 32'hFFFFFFF0;
    // rom_array[5622] = 32'hFFFFFFF0;
    // rom_array[5623] = 32'hFFFFFFF0;
    // rom_array[5624] = 32'hFFFFFFF0;
    // rom_array[5625] = 32'hFFFFFFF0;
    // rom_array[5626] = 32'hFFFFFFF0;
    // rom_array[5627] = 32'hFFFFFFF0;
    // rom_array[5628] = 32'hFFFFFFF0;
    // rom_array[5629] = 32'h000033b9;
    // rom_array[5630] = 32'h000033c1;
    // rom_array[5631] = 32'h000033c9;
    // rom_array[5632] = 32'h000033d1;
    // rom_array[5633] = 32'hFFFFFFF0;
    // rom_array[5634] = 32'hFFFFFFF0;
    // rom_array[5635] = 32'hFFFFFFF0;
    // rom_array[5636] = 32'hFFFFFFF0;
    // rom_array[5637] = 32'h000033d9;
    // rom_array[5638] = 32'h000033e1;
    // rom_array[5639] = 32'h000033e9;
    // rom_array[5640] = 32'h000033f1;
    // rom_array[5641] = 32'h000033f9;
    // rom_array[5642] = 32'h00003401;
    // rom_array[5643] = 32'hFFFFFFF1;
    // rom_array[5644] = 32'hFFFFFFF1;
    // rom_array[5645] = 32'h00003409;
    // rom_array[5646] = 32'h00003411;
    // rom_array[5647] = 32'hFFFFFFF1;
    // rom_array[5648] = 32'hFFFFFFF1;
    // rom_array[5649] = 32'hFFFFFFF0;
    // rom_array[5650] = 32'hFFFFFFF0;
    // rom_array[5651] = 32'hFFFFFFF0;
    // rom_array[5652] = 32'hFFFFFFF0;
    // rom_array[5653] = 32'h00003419;
    // rom_array[5654] = 32'h00003421;
    // rom_array[5655] = 32'hFFFFFFF0;
    // rom_array[5656] = 32'hFFFFFFF0;
    // rom_array[5657] = 32'h00003429;
    // rom_array[5658] = 32'h00003431;
    // rom_array[5659] = 32'hFFFFFFF0;
    // rom_array[5660] = 32'hFFFFFFF0;
    // rom_array[5661] = 32'h00003439;
    // rom_array[5662] = 32'h00003441;
    // rom_array[5663] = 32'hFFFFFFF0;
    // rom_array[5664] = 32'hFFFFFFF0;
    // rom_array[5665] = 32'h00003449;
    // rom_array[5666] = 32'h00003451;
    // rom_array[5667] = 32'hFFFFFFF1;
    // rom_array[5668] = 32'hFFFFFFF1;
    // rom_array[5669] = 32'h00003459;
    // rom_array[5670] = 32'h00003461;
    // rom_array[5671] = 32'hFFFFFFF1;
    // rom_array[5672] = 32'hFFFFFFF1;
    // rom_array[5673] = 32'h00003469;
    // rom_array[5674] = 32'h00003471;
    // rom_array[5675] = 32'hFFFFFFF1;
    // rom_array[5676] = 32'hFFFFFFF1;
    // rom_array[5677] = 32'h00003479;
    // rom_array[5678] = 32'h00003481;
    // rom_array[5679] = 32'hFFFFFFF1;
    // rom_array[5680] = 32'hFFFFFFF1;
    // rom_array[5681] = 32'h00003489;
    // rom_array[5682] = 32'h00003491;
    // rom_array[5683] = 32'hFFFFFFF1;
    // rom_array[5684] = 32'hFFFFFFF1;
    // rom_array[5685] = 32'h00003499;
    // rom_array[5686] = 32'h000034a1;
    // rom_array[5687] = 32'hFFFFFFF1;
    // rom_array[5688] = 32'hFFFFFFF1;
    // rom_array[5689] = 32'h000034a9;
    // rom_array[5690] = 32'h000034b1;
    // rom_array[5691] = 32'hFFFFFFF1;
    // rom_array[5692] = 32'hFFFFFFF1;
    // rom_array[5693] = 32'h000034b9;
    // rom_array[5694] = 32'h000034c1;
    // rom_array[5695] = 32'hFFFFFFF1;
    // rom_array[5696] = 32'hFFFFFFF1;
    // rom_array[5697] = 32'h000034c9;
    // rom_array[5698] = 32'h000034d1;
    // rom_array[5699] = 32'hFFFFFFF0;
    // rom_array[5700] = 32'hFFFFFFF0;
    // rom_array[5701] = 32'h000034d9;
    // rom_array[5702] = 32'h000034e1;
    // rom_array[5703] = 32'hFFFFFFF0;
    // rom_array[5704] = 32'hFFFFFFF0;
    // rom_array[5705] = 32'h000034e9;
    // rom_array[5706] = 32'h000034f1;
    // rom_array[5707] = 32'h000034f9;
    // rom_array[5708] = 32'h00003501;
    // rom_array[5709] = 32'h00003509;
    // rom_array[5710] = 32'h00003511;
    // rom_array[5711] = 32'hFFFFFFF1;
    // rom_array[5712] = 32'hFFFFFFF1;
    // rom_array[5713] = 32'h00003519;
    // rom_array[5714] = 32'h00003521;
    // rom_array[5715] = 32'h00003529;
    // rom_array[5716] = 32'h00003531;
    // rom_array[5717] = 32'hFFFFFFF1;
    // rom_array[5718] = 32'hFFFFFFF1;
    // rom_array[5719] = 32'hFFFFFFF1;
    // rom_array[5720] = 32'hFFFFFFF1;
    // rom_array[5721] = 32'h00003539;
    // rom_array[5722] = 32'h00003541;
    // rom_array[5723] = 32'h00003549;
    // rom_array[5724] = 32'h00003551;
    // rom_array[5725] = 32'hFFFFFFF1;
    // rom_array[5726] = 32'hFFFFFFF1;
    // rom_array[5727] = 32'hFFFFFFF1;
    // rom_array[5728] = 32'hFFFFFFF1;
    // rom_array[5729] = 32'h00003559;
    // rom_array[5730] = 32'h00003561;
    // rom_array[5731] = 32'h00003569;
    // rom_array[5732] = 32'h00003571;
    // rom_array[5733] = 32'hFFFFFFF1;
    // rom_array[5734] = 32'hFFFFFFF1;
    // rom_array[5735] = 32'hFFFFFFF1;
    // rom_array[5736] = 32'hFFFFFFF1;
    // rom_array[5737] = 32'h00003579;
    // rom_array[5738] = 32'h00003581;
    // rom_array[5739] = 32'hFFFFFFF1;
    // rom_array[5740] = 32'hFFFFFFF1;
    // rom_array[5741] = 32'h00003589;
    // rom_array[5742] = 32'h00003591;
    // rom_array[5743] = 32'hFFFFFFF1;
    // rom_array[5744] = 32'hFFFFFFF1;
    // rom_array[5745] = 32'h00003599;
    // rom_array[5746] = 32'h000035a1;
    // rom_array[5747] = 32'h000035a9;
    // rom_array[5748] = 32'h000035b1;
    // rom_array[5749] = 32'h000035b9;
    // rom_array[5750] = 32'h000035c1;
    // rom_array[5751] = 32'hFFFFFFF0;
    // rom_array[5752] = 32'hFFFFFFF0;
    // rom_array[5753] = 32'h000035c9;
    // rom_array[5754] = 32'h000035d1;
    // rom_array[5755] = 32'h000035d9;
    // rom_array[5756] = 32'h000035e1;
    // rom_array[5757] = 32'hFFFFFFF0;
    // rom_array[5758] = 32'hFFFFFFF0;
    // rom_array[5759] = 32'hFFFFFFF0;
    // rom_array[5760] = 32'hFFFFFFF0;
    // rom_array[5761] = 32'h000035e9;
    // rom_array[5762] = 32'h000035f1;
    // rom_array[5763] = 32'h000035f9;
    // rom_array[5764] = 32'h00003601;
    // rom_array[5765] = 32'hFFFFFFF0;
    // rom_array[5766] = 32'hFFFFFFF0;
    // rom_array[5767] = 32'hFFFFFFF0;
    // rom_array[5768] = 32'hFFFFFFF0;
    // rom_array[5769] = 32'h00003609;
    // rom_array[5770] = 32'h00003611;
    // rom_array[5771] = 32'h00003619;
    // rom_array[5772] = 32'h00003621;
    // rom_array[5773] = 32'hFFFFFFF0;
    // rom_array[5774] = 32'hFFFFFFF0;
    // rom_array[5775] = 32'hFFFFFFF0;
    // rom_array[5776] = 32'hFFFFFFF0;
    // rom_array[5777] = 32'h00003629;
    // rom_array[5778] = 32'h00003631;
    // rom_array[5779] = 32'hFFFFFFF1;
    // rom_array[5780] = 32'hFFFFFFF1;
    // rom_array[5781] = 32'h00003639;
    // rom_array[5782] = 32'h00003641;
    // rom_array[5783] = 32'hFFFFFFF1;
    // rom_array[5784] = 32'hFFFFFFF1;
    // rom_array[5785] = 32'h00003649;
    // rom_array[5786] = 32'h00003651;
    // rom_array[5787] = 32'hFFFFFFF1;
    // rom_array[5788] = 32'hFFFFFFF1;
    // rom_array[5789] = 32'h00003659;
    // rom_array[5790] = 32'h00003661;
    // rom_array[5791] = 32'h00003669;
    // rom_array[5792] = 32'h00003671;
    // rom_array[5793] = 32'hFFFFFFF1;
    // rom_array[5794] = 32'hFFFFFFF1;
    // rom_array[5795] = 32'hFFFFFFF1;
    // rom_array[5796] = 32'hFFFFFFF1;
    // rom_array[5797] = 32'h00003679;
    // rom_array[5798] = 32'h00003681;
    // rom_array[5799] = 32'h00003689;
    // rom_array[5800] = 32'h00003691;
    // rom_array[5801] = 32'h00003699;
    // rom_array[5802] = 32'h000036a1;
    // rom_array[5803] = 32'hFFFFFFF0;
    // rom_array[5804] = 32'hFFFFFFF0;
    // rom_array[5805] = 32'h000036a9;
    // rom_array[5806] = 32'h000036b1;
    // rom_array[5807] = 32'hFFFFFFF0;
    // rom_array[5808] = 32'hFFFFFFF0;
    // rom_array[5809] = 32'h000036b9;
    // rom_array[5810] = 32'h000036c1;
    // rom_array[5811] = 32'hFFFFFFF0;
    // rom_array[5812] = 32'hFFFFFFF0;
    // rom_array[5813] = 32'h000036c9;
    // rom_array[5814] = 32'h000036d1;
    // rom_array[5815] = 32'hFFFFFFF0;
    // rom_array[5816] = 32'hFFFFFFF0;
    // rom_array[5817] = 32'h000036d9;
    // rom_array[5818] = 32'h000036e1;
    // rom_array[5819] = 32'h000036e9;
    // rom_array[5820] = 32'h000036f1;
    // rom_array[5821] = 32'h000036f9;
    // rom_array[5822] = 32'h00003701;
    // rom_array[5823] = 32'hFFFFFFF1;
    // rom_array[5824] = 32'hFFFFFFF1;
    // rom_array[5825] = 32'h00003709;
    // rom_array[5826] = 32'h00003711;
    // rom_array[5827] = 32'h00003719;
    // rom_array[5828] = 32'h00003721;
    // rom_array[5829] = 32'hFFFFFFF1;
    // rom_array[5830] = 32'hFFFFFFF1;
    // rom_array[5831] = 32'hFFFFFFF1;
    // rom_array[5832] = 32'hFFFFFFF1;
    // rom_array[5833] = 32'h00003729;
    // rom_array[5834] = 32'h00003731;
    // rom_array[5835] = 32'h00003739;
    // rom_array[5836] = 32'h00003741;
    // rom_array[5837] = 32'hFFFFFFF1;
    // rom_array[5838] = 32'hFFFFFFF1;
    // rom_array[5839] = 32'hFFFFFFF1;
    // rom_array[5840] = 32'hFFFFFFF1;
    // rom_array[5841] = 32'h00003749;
    // rom_array[5842] = 32'h00003751;
    // rom_array[5843] = 32'h00003759;
    // rom_array[5844] = 32'h00003761;
    // rom_array[5845] = 32'hFFFFFFF1;
    // rom_array[5846] = 32'hFFFFFFF1;
    // rom_array[5847] = 32'h00003769;
    // rom_array[5848] = 32'h00003771;
    // rom_array[5849] = 32'h00003779;
    // rom_array[5850] = 32'h00003781;
    // rom_array[5851] = 32'h00003789;
    // rom_array[5852] = 32'h00003791;
    // rom_array[5853] = 32'h00003799;
    // rom_array[5854] = 32'h000037a1;
    // rom_array[5855] = 32'h000037a9;
    // rom_array[5856] = 32'h000037b1;
    // rom_array[5857] = 32'h000037b9;
    // rom_array[5858] = 32'h000037c1;
    // rom_array[5859] = 32'h000037c9;
    // rom_array[5860] = 32'h000037d1;
    // rom_array[5861] = 32'h000037d9;
    // rom_array[5862] = 32'h000037e1;
    // rom_array[5863] = 32'h000037e9;
    // rom_array[5864] = 32'h000037f1;
    // rom_array[5865] = 32'h000037f9;
    // rom_array[5866] = 32'h00003801;
    // rom_array[5867] = 32'hFFFFFFF1;
    // rom_array[5868] = 32'hFFFFFFF1;
    // rom_array[5869] = 32'h00003809;
    // rom_array[5870] = 32'h00003811;
    // rom_array[5871] = 32'hFFFFFFF1;
    // rom_array[5872] = 32'hFFFFFFF1;
    // rom_array[5873] = 32'h00003819;
    // rom_array[5874] = 32'h00003821;
    // rom_array[5875] = 32'h00003829;
    // rom_array[5876] = 32'h00003831;
    // rom_array[5877] = 32'hFFFFFFF0;
    // rom_array[5878] = 32'hFFFFFFF0;
    // rom_array[5879] = 32'hFFFFFFF0;
    // rom_array[5880] = 32'hFFFFFFF0;
    // rom_array[5881] = 32'h00003839;
    // rom_array[5882] = 32'h00003841;
    // rom_array[5883] = 32'h00003849;
    // rom_array[5884] = 32'h00003851;
    // rom_array[5885] = 32'hFFFFFFF0;
    // rom_array[5886] = 32'hFFFFFFF0;
    // rom_array[5887] = 32'hFFFFFFF0;
    // rom_array[5888] = 32'hFFFFFFF0;
    // rom_array[5889] = 32'hFFFFFFF0;
    // rom_array[5890] = 32'hFFFFFFF0;
    // rom_array[5891] = 32'h00003859;
    // rom_array[5892] = 32'h00003861;
    // rom_array[5893] = 32'hFFFFFFF0;
    // rom_array[5894] = 32'hFFFFFFF0;
    // rom_array[5895] = 32'h00003869;
    // rom_array[5896] = 32'h00003871;
    // rom_array[5897] = 32'h00003879;
    // rom_array[5898] = 32'h00003881;
    // rom_array[5899] = 32'h00003889;
    // rom_array[5900] = 32'h00003891;
    // rom_array[5901] = 32'hFFFFFFF0;
    // rom_array[5902] = 32'hFFFFFFF0;
    // rom_array[5903] = 32'hFFFFFFF0;
    // rom_array[5904] = 32'hFFFFFFF0;
    // rom_array[5905] = 32'h00003899;
    // rom_array[5906] = 32'h000038a1;
    // rom_array[5907] = 32'h000038a9;
    // rom_array[5908] = 32'h000038b1;
    // rom_array[5909] = 32'hFFFFFFF0;
    // rom_array[5910] = 32'hFFFFFFF0;
    // rom_array[5911] = 32'h000038b9;
    // rom_array[5912] = 32'h000038c1;
    // rom_array[5913] = 32'h000038c9;
    // rom_array[5914] = 32'h000038d1;
    // rom_array[5915] = 32'h000038d9;
    // rom_array[5916] = 32'h000038e1;
    // rom_array[5917] = 32'hFFFFFFF0;
    // rom_array[5918] = 32'hFFFFFFF0;
    // rom_array[5919] = 32'hFFFFFFF0;
    // rom_array[5920] = 32'hFFFFFFF0;
    // rom_array[5921] = 32'h000038e9;
    // rom_array[5922] = 32'h000038f1;
    // rom_array[5923] = 32'h000038f9;
    // rom_array[5924] = 32'h00003901;
    // rom_array[5925] = 32'hFFFFFFF0;
    // rom_array[5926] = 32'hFFFFFFF0;
    // rom_array[5927] = 32'hFFFFFFF0;
    // rom_array[5928] = 32'hFFFFFFF0;
    // rom_array[5929] = 32'hFFFFFFF0;
    // rom_array[5930] = 32'hFFFFFFF0;
    // rom_array[5931] = 32'h00003909;
    // rom_array[5932] = 32'h00003911;
    // rom_array[5933] = 32'hFFFFFFF0;
    // rom_array[5934] = 32'hFFFFFFF0;
    // rom_array[5935] = 32'h00003919;
    // rom_array[5936] = 32'h00003921;
    // rom_array[5937] = 32'hFFFFFFF0;
    // rom_array[5938] = 32'hFFFFFFF0;
    // rom_array[5939] = 32'h00003929;
    // rom_array[5940] = 32'h00003931;
    // rom_array[5941] = 32'hFFFFFFF0;
    // rom_array[5942] = 32'hFFFFFFF0;
    // rom_array[5943] = 32'h00003939;
    // rom_array[5944] = 32'h00003941;
    // rom_array[5945] = 32'hFFFFFFF0;
    // rom_array[5946] = 32'hFFFFFFF0;
    // rom_array[5947] = 32'hFFFFFFF0;
    // rom_array[5948] = 32'hFFFFFFF0;
    // rom_array[5949] = 32'hFFFFFFF1;
    // rom_array[5950] = 32'hFFFFFFF1;
    // rom_array[5951] = 32'hFFFFFFF1;
    // rom_array[5952] = 32'hFFFFFFF1;
    // rom_array[5953] = 32'hFFFFFFF0;
    // rom_array[5954] = 32'hFFFFFFF0;
    // rom_array[5955] = 32'hFFFFFFF0;
    // rom_array[5956] = 32'hFFFFFFF0;
    // rom_array[5957] = 32'h00003949;
    // rom_array[5958] = 32'h00003951;
    // rom_array[5959] = 32'hFFFFFFF0;
    // rom_array[5960] = 32'hFFFFFFF0;
    // rom_array[5961] = 32'hFFFFFFF0;
    // rom_array[5962] = 32'hFFFFFFF0;
    // rom_array[5963] = 32'h00003959;
    // rom_array[5964] = 32'h00003961;
    // rom_array[5965] = 32'hFFFFFFF0;
    // rom_array[5966] = 32'hFFFFFFF0;
    // rom_array[5967] = 32'h00003969;
    // rom_array[5968] = 32'h00003971;
    // rom_array[5969] = 32'hFFFFFFF0;
    // rom_array[5970] = 32'hFFFFFFF0;
    // rom_array[5971] = 32'h00003979;
    // rom_array[5972] = 32'h00003981;
    // rom_array[5973] = 32'hFFFFFFF0;
    // rom_array[5974] = 32'hFFFFFFF0;
    // rom_array[5975] = 32'h00003989;
    // rom_array[5976] = 32'h00003991;
    // rom_array[5977] = 32'h00003999;
    // rom_array[5978] = 32'h000039a1;
    // rom_array[5979] = 32'h000039a9;
    // rom_array[5980] = 32'h000039b1;
    // rom_array[5981] = 32'hFFFFFFF1;
    // rom_array[5982] = 32'hFFFFFFF1;
    // rom_array[5983] = 32'hFFFFFFF1;
    // rom_array[5984] = 32'hFFFFFFF1;
    // rom_array[5985] = 32'h000039b9;
    // rom_array[5986] = 32'h000039c1;
    // rom_array[5987] = 32'h000039c9;
    // rom_array[5988] = 32'h000039d1;
    // rom_array[5989] = 32'h000039d9;
    // rom_array[5990] = 32'h000039e1;
    // rom_array[5991] = 32'hFFFFFFF1;
    // rom_array[5992] = 32'hFFFFFFF1;
    // rom_array[5993] = 32'h000039e9;
    // rom_array[5994] = 32'h000039f1;
    // rom_array[5995] = 32'h000039f9;
    // rom_array[5996] = 32'h00003a01;
    // rom_array[5997] = 32'hFFFFFFF0;
    // rom_array[5998] = 32'hFFFFFFF0;
    // rom_array[5999] = 32'hFFFFFFF0;
    // rom_array[6000] = 32'hFFFFFFF0;
    // rom_array[6001] = 32'h00003a09;
    // rom_array[6002] = 32'h00003a11;
    // rom_array[6003] = 32'h00003a19;
    // rom_array[6004] = 32'h00003a21;
    // rom_array[6005] = 32'h00003a29;
    // rom_array[6006] = 32'h00003a31;
    // rom_array[6007] = 32'hFFFFFFF0;
    // rom_array[6008] = 32'hFFFFFFF0;
    // rom_array[6009] = 32'hFFFFFFF0;
    // rom_array[6010] = 32'hFFFFFFF0;
    // rom_array[6011] = 32'h00003a39;
    // rom_array[6012] = 32'h00003a41;
    // rom_array[6013] = 32'hFFFFFFF0;
    // rom_array[6014] = 32'hFFFFFFF0;
    // rom_array[6015] = 32'h00003a49;
    // rom_array[6016] = 32'h00003a51;
    // rom_array[6017] = 32'hFFFFFFF0;
    // rom_array[6018] = 32'hFFFFFFF0;
    // rom_array[6019] = 32'h00003a59;
    // rom_array[6020] = 32'h00003a61;
    // rom_array[6021] = 32'hFFFFFFF0;
    // rom_array[6022] = 32'hFFFFFFF0;
    // rom_array[6023] = 32'h00003a69;
    // rom_array[6024] = 32'h00003a71;
    // rom_array[6025] = 32'h00003a79;
    // rom_array[6026] = 32'h00003a81;
    // rom_array[6027] = 32'h00003a89;
    // rom_array[6028] = 32'h00003a91;
    // rom_array[6029] = 32'h00003a99;
    // rom_array[6030] = 32'h00003aa1;
    // rom_array[6031] = 32'hFFFFFFF1;
    // rom_array[6032] = 32'hFFFFFFF1;
    // rom_array[6033] = 32'h00003aa9;
    // rom_array[6034] = 32'h00003ab1;
    // rom_array[6035] = 32'h00003ab9;
    // rom_array[6036] = 32'h00003ac1;
    // rom_array[6037] = 32'hFFFFFFF1;
    // rom_array[6038] = 32'hFFFFFFF1;
    // rom_array[6039] = 32'hFFFFFFF1;
    // rom_array[6040] = 32'hFFFFFFF1;
    // rom_array[6041] = 32'h00003ac9;
    // rom_array[6042] = 32'h00003ad1;
    // rom_array[6043] = 32'hFFFFFFF1;
    // rom_array[6044] = 32'hFFFFFFF1;
    // rom_array[6045] = 32'h00003ad9;
    // rom_array[6046] = 32'h00003ae1;
    // rom_array[6047] = 32'hFFFFFFF1;
    // rom_array[6048] = 32'hFFFFFFF1;
    // rom_array[6049] = 32'h00003ae9;
    // rom_array[6050] = 32'h00003af1;
    // rom_array[6051] = 32'h00003af9;
    // rom_array[6052] = 32'h00003b01;
    // rom_array[6053] = 32'hFFFFFFF0;
    // rom_array[6054] = 32'hFFFFFFF0;
    // rom_array[6055] = 32'hFFFFFFF0;
    // rom_array[6056] = 32'hFFFFFFF0;
    // rom_array[6057] = 32'h00003b09;
    // rom_array[6058] = 32'h00003b11;
    // rom_array[6059] = 32'h00003b19;
    // rom_array[6060] = 32'h00003b21;
    // rom_array[6061] = 32'hFFFFFFF0;
    // rom_array[6062] = 32'hFFFFFFF0;
    // rom_array[6063] = 32'hFFFFFFF0;
    // rom_array[6064] = 32'hFFFFFFF0;
    // rom_array[6065] = 32'h00003b29;
    // rom_array[6066] = 32'h00003b31;
    // rom_array[6067] = 32'h00003b39;
    // rom_array[6068] = 32'h00003b41;
    // rom_array[6069] = 32'hFFFFFFF1;
    // rom_array[6070] = 32'hFFFFFFF1;
    // rom_array[6071] = 32'hFFFFFFF1;
    // rom_array[6072] = 32'hFFFFFFF1;
    // rom_array[6073] = 32'h00003b49;
    // rom_array[6074] = 32'h00003b51;
    // rom_array[6075] = 32'h00003b59;
    // rom_array[6076] = 32'h00003b61;
    // rom_array[6077] = 32'hFFFFFFF1;
    // rom_array[6078] = 32'hFFFFFFF1;
    // rom_array[6079] = 32'h00003b69;
    // rom_array[6080] = 32'h00003b71;
    // rom_array[6081] = 32'hFFFFFFF0;
    // rom_array[6082] = 32'hFFFFFFF0;
    // rom_array[6083] = 32'h00003b79;
    // rom_array[6084] = 32'h00003b81;
    // rom_array[6085] = 32'hFFFFFFF0;
    // rom_array[6086] = 32'hFFFFFFF0;
    // rom_array[6087] = 32'h00003b89;
    // rom_array[6088] = 32'h00003b91;
    // rom_array[6089] = 32'h00003b99;
    // rom_array[6090] = 32'h00003ba1;
    // rom_array[6091] = 32'h00003ba9;
    // rom_array[6092] = 32'h00003bb1;
    // rom_array[6093] = 32'hFFFFFFF1;
    // rom_array[6094] = 32'hFFFFFFF1;
    // rom_array[6095] = 32'hFFFFFFF1;
    // rom_array[6096] = 32'hFFFFFFF1;
    // rom_array[6097] = 32'h00003bb9;
    // rom_array[6098] = 32'h00003bc1;
    // rom_array[6099] = 32'h00003bc9;
    // rom_array[6100] = 32'h00003bd1;
    // rom_array[6101] = 32'hFFFFFFF1;
    // rom_array[6102] = 32'hFFFFFFF1;
    // rom_array[6103] = 32'hFFFFFFF1;
    // rom_array[6104] = 32'hFFFFFFF1;
    // rom_array[6105] = 32'hFFFFFFF1;
    // rom_array[6106] = 32'hFFFFFFF1;
    // rom_array[6107] = 32'hFFFFFFF1;
    // rom_array[6108] = 32'hFFFFFFF1;
    // rom_array[6109] = 32'h00003bd9;
    // rom_array[6110] = 32'h00003be1;
    // rom_array[6111] = 32'h00003be9;
    // rom_array[6112] = 32'h00003bf1;
    // rom_array[6113] = 32'hFFFFFFF1;
    // rom_array[6114] = 32'hFFFFFFF1;
    // rom_array[6115] = 32'hFFFFFFF1;
    // rom_array[6116] = 32'hFFFFFFF1;
    // rom_array[6117] = 32'h00003bf9;
    // rom_array[6118] = 32'h00003c01;
    // rom_array[6119] = 32'h00003c09;
    // rom_array[6120] = 32'h00003c11;
    // rom_array[6121] = 32'h00003c19;
    // rom_array[6122] = 32'h00003c21;
    // rom_array[6123] = 32'h00003c29;
    // rom_array[6124] = 32'h00003c31;
    // rom_array[6125] = 32'hFFFFFFF0;
    // rom_array[6126] = 32'hFFFFFFF0;
    // rom_array[6127] = 32'hFFFFFFF0;
    // rom_array[6128] = 32'hFFFFFFF0;
    // rom_array[6129] = 32'h00003c39;
    // rom_array[6130] = 32'h00003c41;
    // rom_array[6131] = 32'h00003c49;
    // rom_array[6132] = 32'h00003c51;
    // rom_array[6133] = 32'hFFFFFFF0;
    // rom_array[6134] = 32'hFFFFFFF0;
    // rom_array[6135] = 32'hFFFFFFF0;
    // rom_array[6136] = 32'hFFFFFFF0;
    // rom_array[6137] = 32'h00003c59;
    // rom_array[6138] = 32'h00003c61;
    // rom_array[6139] = 32'h00003c69;
    // rom_array[6140] = 32'h00003c71;
    // rom_array[6141] = 32'hFFFFFFF0;
    // rom_array[6142] = 32'hFFFFFFF0;
    // rom_array[6143] = 32'hFFFFFFF0;
    // rom_array[6144] = 32'hFFFFFFF0;
    // rom_array[6145] = 32'h00003c79;
    // rom_array[6146] = 32'h00003c81;
    // rom_array[6147] = 32'h00003c89;
    // rom_array[6148] = 32'h00003c91;
    // rom_array[6149] = 32'hFFFFFFF0;
    // rom_array[6150] = 32'hFFFFFFF0;
    // rom_array[6151] = 32'hFFFFFFF0;
    // rom_array[6152] = 32'hFFFFFFF0;
    // rom_array[6153] = 32'h00003c99;
    // rom_array[6154] = 32'h00003ca1;
    // rom_array[6155] = 32'h00003ca9;
    // rom_array[6156] = 32'h00003cb1;
    // rom_array[6157] = 32'h00003cb9;
    // rom_array[6158] = 32'h00003cc1;
    // rom_array[6159] = 32'hFFFFFFF1;
    // rom_array[6160] = 32'hFFFFFFF1;
    // rom_array[6161] = 32'h00003cc9;
    // rom_array[6162] = 32'h00003cd1;
    // rom_array[6163] = 32'h00003cd9;
    // rom_array[6164] = 32'h00003ce1;
    // rom_array[6165] = 32'hFFFFFFF1;
    // rom_array[6166] = 32'hFFFFFFF1;
    // rom_array[6167] = 32'hFFFFFFF1;
    // rom_array[6168] = 32'hFFFFFFF1;
    // rom_array[6169] = 32'h00003ce9;
    // rom_array[6170] = 32'h00003cf1;
    // rom_array[6171] = 32'hFFFFFFF1;
    // rom_array[6172] = 32'hFFFFFFF1;
    // rom_array[6173] = 32'h00003cf9;
    // rom_array[6174] = 32'h00003d01;
    // rom_array[6175] = 32'hFFFFFFF1;
    // rom_array[6176] = 32'hFFFFFFF1;
    // rom_array[6177] = 32'h00003d09;
    // rom_array[6178] = 32'h00003d11;
    // rom_array[6179] = 32'h00003d19;
    // rom_array[6180] = 32'h00003d21;
    // rom_array[6181] = 32'hFFFFFFF0;
    // rom_array[6182] = 32'hFFFFFFF0;
    // rom_array[6183] = 32'hFFFFFFF0;
    // rom_array[6184] = 32'hFFFFFFF0;
    // rom_array[6185] = 32'h00003d29;
    // rom_array[6186] = 32'h00003d31;
    // rom_array[6187] = 32'h00003d39;
    // rom_array[6188] = 32'h00003d41;
    // rom_array[6189] = 32'hFFFFFFF0;
    // rom_array[6190] = 32'hFFFFFFF0;
    // rom_array[6191] = 32'hFFFFFFF0;
    // rom_array[6192] = 32'hFFFFFFF0;
    // rom_array[6193] = 32'h00003d49;
    // rom_array[6194] = 32'h00003d51;
    // rom_array[6195] = 32'h00003d59;
    // rom_array[6196] = 32'h00003d61;
    // rom_array[6197] = 32'hFFFFFFF1;
    // rom_array[6198] = 32'hFFFFFFF1;
    // rom_array[6199] = 32'hFFFFFFF1;
    // rom_array[6200] = 32'hFFFFFFF1;
    // rom_array[6201] = 32'h00003d69;
    // rom_array[6202] = 32'h00003d71;
    // rom_array[6203] = 32'h00003d79;
    // rom_array[6204] = 32'h00003d81;
    // rom_array[6205] = 32'hFFFFFFF1;
    // rom_array[6206] = 32'hFFFFFFF1;
    // rom_array[6207] = 32'hFFFFFFF1;
    // rom_array[6208] = 32'hFFFFFFF1;
    // rom_array[6209] = 32'h00003d89;
    // rom_array[6210] = 32'h00003d91;
    // rom_array[6211] = 32'h00003d99;
    // rom_array[6212] = 32'h00003da1;
    // rom_array[6213] = 32'hFFFFFFF1;
    // rom_array[6214] = 32'hFFFFFFF1;
    // rom_array[6215] = 32'hFFFFFFF1;
    // rom_array[6216] = 32'hFFFFFFF1;
    // rom_array[6217] = 32'h00003da9;
    // rom_array[6218] = 32'h00003db1;
    // rom_array[6219] = 32'h00003db9;
    // rom_array[6220] = 32'h00003dc1;
    // rom_array[6221] = 32'hFFFFFFF1;
    // rom_array[6222] = 32'hFFFFFFF1;
    // rom_array[6223] = 32'hFFFFFFF1;
    // rom_array[6224] = 32'hFFFFFFF1;
    // rom_array[6225] = 32'h00003dc9;
    // rom_array[6226] = 32'h00003dd1;
    // rom_array[6227] = 32'h00003dd9;
    // rom_array[6228] = 32'h00003de1;
    // rom_array[6229] = 32'hFFFFFFF0;
    // rom_array[6230] = 32'hFFFFFFF0;
    // rom_array[6231] = 32'hFFFFFFF0;
    // rom_array[6232] = 32'hFFFFFFF0;
    // rom_array[6233] = 32'h00003de9;
    // rom_array[6234] = 32'h00003df1;
    // rom_array[6235] = 32'h00003df9;
    // rom_array[6236] = 32'h00003e01;
    // rom_array[6237] = 32'hFFFFFFF0;
    // rom_array[6238] = 32'hFFFFFFF0;
    // rom_array[6239] = 32'hFFFFFFF0;
    // rom_array[6240] = 32'hFFFFFFF0;
    // rom_array[6241] = 32'h00003e09;
    // rom_array[6242] = 32'h00003e11;
    // rom_array[6243] = 32'h00003e19;
    // rom_array[6244] = 32'h00003e21;
    // rom_array[6245] = 32'h00003e29;
    // rom_array[6246] = 32'h00003e31;
    // rom_array[6247] = 32'hFFFFFFF1;
    // rom_array[6248] = 32'hFFFFFFF1;
    // rom_array[6249] = 32'h00003e39;
    // rom_array[6250] = 32'h00003e41;
    // rom_array[6251] = 32'h00003e49;
    // rom_array[6252] = 32'h00003e51;
    // rom_array[6253] = 32'hFFFFFFF1;
    // rom_array[6254] = 32'hFFFFFFF1;
    // rom_array[6255] = 32'hFFFFFFF1;
    // rom_array[6256] = 32'hFFFFFFF1;
    // rom_array[6257] = 32'h00003e59;
    // rom_array[6258] = 32'h00003e61;
    // rom_array[6259] = 32'hFFFFFFF1;
    // rom_array[6260] = 32'hFFFFFFF1;
    // rom_array[6261] = 32'h00003e69;
    // rom_array[6262] = 32'h00003e71;
    // rom_array[6263] = 32'hFFFFFFF1;
    // rom_array[6264] = 32'hFFFFFFF1;
    // rom_array[6265] = 32'h00003e79;
    // rom_array[6266] = 32'h00003e81;
    // rom_array[6267] = 32'hFFFFFFF1;
    // rom_array[6268] = 32'hFFFFFFF1;
    // rom_array[6269] = 32'h00003e89;
    // rom_array[6270] = 32'h00003e91;
    // rom_array[6271] = 32'hFFFFFFF1;
    // rom_array[6272] = 32'hFFFFFFF1;
    // rom_array[6273] = 32'h00003e99;
    // rom_array[6274] = 32'h00003ea1;
    // rom_array[6275] = 32'hFFFFFFF1;
    // rom_array[6276] = 32'hFFFFFFF1;
    // rom_array[6277] = 32'h00003ea9;
    // rom_array[6278] = 32'h00003eb1;
    // rom_array[6279] = 32'hFFFFFFF1;
    // rom_array[6280] = 32'hFFFFFFF1;
    // rom_array[6281] = 32'hFFFFFFF0;
    // rom_array[6282] = 32'hFFFFFFF0;
    // rom_array[6283] = 32'hFFFFFFF0;
    // rom_array[6284] = 32'hFFFFFFF0;
    // rom_array[6285] = 32'hFFFFFFF0;
    // rom_array[6286] = 32'hFFFFFFF0;
    // rom_array[6287] = 32'h00003eb9;
    // rom_array[6288] = 32'h00003ec1;
    // rom_array[6289] = 32'h00003ec9;
    // rom_array[6290] = 32'h00003ed1;
    // rom_array[6291] = 32'h00003ed9;
    // rom_array[6292] = 32'h00003ee1;
    // rom_array[6293] = 32'hFFFFFFF0;
    // rom_array[6294] = 32'hFFFFFFF0;
    // rom_array[6295] = 32'hFFFFFFF0;
    // rom_array[6296] = 32'hFFFFFFF0;
    // rom_array[6297] = 32'h00003ee9;
    // rom_array[6298] = 32'h00003ef1;
    // rom_array[6299] = 32'h00003ef9;
    // rom_array[6300] = 32'h00003f01;
    // rom_array[6301] = 32'hFFFFFFF0;
    // rom_array[6302] = 32'hFFFFFFF0;
    // rom_array[6303] = 32'h00003f09;
    // rom_array[6304] = 32'h00003f11;
    // rom_array[6305] = 32'hFFFFFFF0;
    // rom_array[6306] = 32'hFFFFFFF0;
    // rom_array[6307] = 32'h00003f19;
    // rom_array[6308] = 32'h00003f21;
    // rom_array[6309] = 32'hFFFFFFF0;
    // rom_array[6310] = 32'hFFFFFFF0;
    // rom_array[6311] = 32'h00003f29;
    // rom_array[6312] = 32'h00003f31;
    // rom_array[6313] = 32'h00003f39;
    // rom_array[6314] = 32'h00003f41;
    // rom_array[6315] = 32'h00003f49;
    // rom_array[6316] = 32'h00003f51;
    // rom_array[6317] = 32'h00003f59;
    // rom_array[6318] = 32'h00003f61;
    // rom_array[6319] = 32'hFFFFFFF1;
    // rom_array[6320] = 32'hFFFFFFF1;
    // rom_array[6321] = 32'h00003f69;
    // rom_array[6322] = 32'h00003f71;
    // rom_array[6323] = 32'h00003f79;
    // rom_array[6324] = 32'h00003f81;
    // rom_array[6325] = 32'hFFFFFFF1;
    // rom_array[6326] = 32'hFFFFFFF1;
    // rom_array[6327] = 32'hFFFFFFF1;
    // rom_array[6328] = 32'hFFFFFFF1;
    // rom_array[6329] = 32'h00003f89;
    // rom_array[6330] = 32'h00003f91;
    // rom_array[6331] = 32'hFFFFFFF1;
    // rom_array[6332] = 32'hFFFFFFF1;
    // rom_array[6333] = 32'h00003f99;
    // rom_array[6334] = 32'h00003fa1;
    // rom_array[6335] = 32'hFFFFFFF1;
    // rom_array[6336] = 32'hFFFFFFF1;
    // rom_array[6337] = 32'h00003fa9;
    // rom_array[6338] = 32'h00003fb1;
    // rom_array[6339] = 32'h00003fb9;
    // rom_array[6340] = 32'h00003fc1;
    // rom_array[6341] = 32'h00003fc9;
    // rom_array[6342] = 32'h00003fd1;
    // rom_array[6343] = 32'hFFFFFFF1;
    // rom_array[6344] = 32'hFFFFFFF1;
    // rom_array[6345] = 32'h00003fd9;
    // rom_array[6346] = 32'h00003fe1;
    // rom_array[6347] = 32'h00003fe9;
    // rom_array[6348] = 32'h00003ff1;
    // rom_array[6349] = 32'hFFFFFFF1;
    // rom_array[6350] = 32'hFFFFFFF1;
    // rom_array[6351] = 32'hFFFFFFF1;
    // rom_array[6352] = 32'hFFFFFFF1;
    // rom_array[6353] = 32'h00003ff9;
    // rom_array[6354] = 32'h00004001;
    // rom_array[6355] = 32'h00004009;
    // rom_array[6356] = 32'h00004011;
    // rom_array[6357] = 32'hFFFFFFF1;
    // rom_array[6358] = 32'hFFFFFFF1;
    // rom_array[6359] = 32'hFFFFFFF1;
    // rom_array[6360] = 32'hFFFFFFF1;
    // rom_array[6361] = 32'h00004019;
    // rom_array[6362] = 32'h00004021;
    // rom_array[6363] = 32'h00004029;
    // rom_array[6364] = 32'h00004031;
    // rom_array[6365] = 32'hFFFFFFF1;
    // rom_array[6366] = 32'hFFFFFFF1;
    // rom_array[6367] = 32'hFFFFFFF1;
    // rom_array[6368] = 32'hFFFFFFF1;
    // rom_array[6369] = 32'h00004039;
    // rom_array[6370] = 32'h00004041;
    // rom_array[6371] = 32'h00004049;
    // rom_array[6372] = 32'h00004051;
    // rom_array[6373] = 32'hFFFFFFF1;
    // rom_array[6374] = 32'hFFFFFFF1;
    // rom_array[6375] = 32'hFFFFFFF1;
    // rom_array[6376] = 32'hFFFFFFF1;
    // rom_array[6377] = 32'h00004059;
    // rom_array[6378] = 32'h00004061;
    // rom_array[6379] = 32'h00004069;
    // rom_array[6380] = 32'h00004071;
    // rom_array[6381] = 32'hFFFFFFF1;
    // rom_array[6382] = 32'hFFFFFFF1;
    // rom_array[6383] = 32'hFFFFFFF1;
    // rom_array[6384] = 32'hFFFFFFF1;
    // rom_array[6385] = 32'h00004079;
    // rom_array[6386] = 32'h00004081;
    // rom_array[6387] = 32'h00004089;
    // rom_array[6388] = 32'h00004091;
    // rom_array[6389] = 32'h00004099;
    // rom_array[6390] = 32'h000040a1;
    // rom_array[6391] = 32'hFFFFFFF0;
    // rom_array[6392] = 32'hFFFFFFF0;
    // rom_array[6393] = 32'h000040a9;
    // rom_array[6394] = 32'h000040b1;
    // rom_array[6395] = 32'h000040b9;
    // rom_array[6396] = 32'h000040c1;
    // rom_array[6397] = 32'hFFFFFFF0;
    // rom_array[6398] = 32'hFFFFFFF0;
    // rom_array[6399] = 32'hFFFFFFF0;
    // rom_array[6400] = 32'hFFFFFFF0;
    // rom_array[6401] = 32'h000040c9;
    // rom_array[6402] = 32'h000040d1;
    // rom_array[6403] = 32'h000040d9;
    // rom_array[6404] = 32'h000040e1;
    // rom_array[6405] = 32'hFFFFFFF0;
    // rom_array[6406] = 32'hFFFFFFF0;
    // rom_array[6407] = 32'h000040e9;
    // rom_array[6408] = 32'h000040f1;
    // rom_array[6409] = 32'h000040f9;
    // rom_array[6410] = 32'h00004101;
    // rom_array[6411] = 32'h00004109;
    // rom_array[6412] = 32'h00004111;
    // rom_array[6413] = 32'hFFFFFFF1;
    // rom_array[6414] = 32'hFFFFFFF1;
    // rom_array[6415] = 32'hFFFFFFF1;
    // rom_array[6416] = 32'hFFFFFFF1;
    // rom_array[6417] = 32'h00004119;
    // rom_array[6418] = 32'h00004121;
    // rom_array[6419] = 32'hFFFFFFF1;
    // rom_array[6420] = 32'hFFFFFFF1;
    // rom_array[6421] = 32'h00004129;
    // rom_array[6422] = 32'h00004131;
    // rom_array[6423] = 32'hFFFFFFF1;
    // rom_array[6424] = 32'hFFFFFFF1;
    // rom_array[6425] = 32'h00004139;
    // rom_array[6426] = 32'h00004141;
    // rom_array[6427] = 32'hFFFFFFF1;
    // rom_array[6428] = 32'hFFFFFFF1;
    // rom_array[6429] = 32'h00004149;
    // rom_array[6430] = 32'h00004151;
    // rom_array[6431] = 32'hFFFFFFF1;
    // rom_array[6432] = 32'hFFFFFFF1;
    // rom_array[6433] = 32'h00004159;
    // rom_array[6434] = 32'h00004161;
    // rom_array[6435] = 32'hFFFFFFF1;
    // rom_array[6436] = 32'hFFFFFFF1;
    // rom_array[6437] = 32'h00004169;
    // rom_array[6438] = 32'h00004171;
    // rom_array[6439] = 32'hFFFFFFF1;
    // rom_array[6440] = 32'hFFFFFFF1;
    // rom_array[6441] = 32'h00004179;
    // rom_array[6442] = 32'h00004181;
    // rom_array[6443] = 32'hFFFFFFF1;
    // rom_array[6444] = 32'hFFFFFFF1;
    // rom_array[6445] = 32'h00004189;
    // rom_array[6446] = 32'h00004191;
    // rom_array[6447] = 32'hFFFFFFF1;
    // rom_array[6448] = 32'hFFFFFFF1;
    // rom_array[6449] = 32'h00004199;
    // rom_array[6450] = 32'h000041a1;
    // rom_array[6451] = 32'hFFFFFFF0;
    // rom_array[6452] = 32'hFFFFFFF0;
    // rom_array[6453] = 32'h000041a9;
    // rom_array[6454] = 32'h000041b1;
    // rom_array[6455] = 32'hFFFFFFF0;
    // rom_array[6456] = 32'hFFFFFFF0;
    // rom_array[6457] = 32'h000041b9;
    // rom_array[6458] = 32'h000041c1;
    // rom_array[6459] = 32'hFFFFFFF0;
    // rom_array[6460] = 32'hFFFFFFF0;
    // rom_array[6461] = 32'h000041c9;
    // rom_array[6462] = 32'h000041d1;
    // rom_array[6463] = 32'hFFFFFFF0;
    // rom_array[6464] = 32'hFFFFFFF0;
    // rom_array[6465] = 32'hFFFFFFF0;
    // rom_array[6466] = 32'hFFFFFFF0;
    // rom_array[6467] = 32'h000041d9;
    // rom_array[6468] = 32'h000041e1;
    // rom_array[6469] = 32'hFFFFFFF0;
    // rom_array[6470] = 32'hFFFFFFF0;
    // rom_array[6471] = 32'h000041e9;
    // rom_array[6472] = 32'h000041f1;
    // rom_array[6473] = 32'hFFFFFFF0;
    // rom_array[6474] = 32'hFFFFFFF0;
    // rom_array[6475] = 32'h000041f9;
    // rom_array[6476] = 32'h00004201;
    // rom_array[6477] = 32'hFFFFFFF0;
    // rom_array[6478] = 32'hFFFFFFF0;
    // rom_array[6479] = 32'h00004209;
    // rom_array[6480] = 32'h00004211;
    // rom_array[6481] = 32'h00004219;
    // rom_array[6482] = 32'h00004221;
    // rom_array[6483] = 32'hFFFFFFF0;
    // rom_array[6484] = 32'hFFFFFFF0;
    // rom_array[6485] = 32'h00004229;
    // rom_array[6486] = 32'h00004231;
    // rom_array[6487] = 32'hFFFFFFF0;
    // rom_array[6488] = 32'hFFFFFFF0;
    // rom_array[6489] = 32'h00004239;
    // rom_array[6490] = 32'h00004241;
    // rom_array[6491] = 32'hFFFFFFF0;
    // rom_array[6492] = 32'hFFFFFFF0;
    // rom_array[6493] = 32'h00004249;
    // rom_array[6494] = 32'h00004251;
    // rom_array[6495] = 32'hFFFFFFF0;
    // rom_array[6496] = 32'hFFFFFFF0;
    // rom_array[6497] = 32'hFFFFFFF0;
    // rom_array[6498] = 32'hFFFFFFF0;
    // rom_array[6499] = 32'h00004259;
    // rom_array[6500] = 32'h00004261;
    // rom_array[6501] = 32'hFFFFFFF0;
    // rom_array[6502] = 32'hFFFFFFF0;
    // rom_array[6503] = 32'h00004269;
    // rom_array[6504] = 32'h00004271;
    // rom_array[6505] = 32'hFFFFFFF0;
    // rom_array[6506] = 32'hFFFFFFF0;
    // rom_array[6507] = 32'h00004279;
    // rom_array[6508] = 32'h00004281;
    // rom_array[6509] = 32'hFFFFFFF0;
    // rom_array[6510] = 32'hFFFFFFF0;
    // rom_array[6511] = 32'h00004289;
    // rom_array[6512] = 32'h00004291;
    // rom_array[6513] = 32'hFFFFFFF0;
    // rom_array[6514] = 32'hFFFFFFF0;
    // rom_array[6515] = 32'hFFFFFFF0;
    // rom_array[6516] = 32'hFFFFFFF0;
    // rom_array[6517] = 32'h00004299;
    // rom_array[6518] = 32'h000042a1;
    // rom_array[6519] = 32'h000042a9;
    // rom_array[6520] = 32'h000042b1;
    // rom_array[6521] = 32'hFFFFFFF0;
    // rom_array[6522] = 32'hFFFFFFF0;
    // rom_array[6523] = 32'hFFFFFFF0;
    // rom_array[6524] = 32'hFFFFFFF0;
    // rom_array[6525] = 32'h000042b9;
    // rom_array[6526] = 32'h000042c1;
    // rom_array[6527] = 32'h000042c9;
    // rom_array[6528] = 32'h000042d1;
    // rom_array[6529] = 32'h000042d9;
    // rom_array[6530] = 32'h000042e1;
    // rom_array[6531] = 32'hFFFFFFF1;
    // rom_array[6532] = 32'hFFFFFFF1;
    // rom_array[6533] = 32'h000042e9;
    // rom_array[6534] = 32'h000042f1;
    // rom_array[6535] = 32'hFFFFFFF1;
    // rom_array[6536] = 32'hFFFFFFF1;
    // rom_array[6537] = 32'hFFFFFFF0;
    // rom_array[6538] = 32'hFFFFFFF0;
    // rom_array[6539] = 32'hFFFFFFF0;
    // rom_array[6540] = 32'hFFFFFFF0;
    // rom_array[6541] = 32'h000042f9;
    // rom_array[6542] = 32'h00004301;
    // rom_array[6543] = 32'hFFFFFFF0;
    // rom_array[6544] = 32'hFFFFFFF0;
    // rom_array[6545] = 32'h00004309;
    // rom_array[6546] = 32'h00004311;
    // rom_array[6547] = 32'hFFFFFFF0;
    // rom_array[6548] = 32'hFFFFFFF0;
    // rom_array[6549] = 32'h00004319;
    // rom_array[6550] = 32'h00004321;
    // rom_array[6551] = 32'hFFFFFFF0;
    // rom_array[6552] = 32'hFFFFFFF0;
    // rom_array[6553] = 32'h00004329;
    // rom_array[6554] = 32'h00004331;
    // rom_array[6555] = 32'hFFFFFFF1;
    // rom_array[6556] = 32'hFFFFFFF1;
    // rom_array[6557] = 32'h00004339;
    // rom_array[6558] = 32'h00004341;
    // rom_array[6559] = 32'hFFFFFFF1;
    // rom_array[6560] = 32'hFFFFFFF1;
    // rom_array[6561] = 32'h00004349;
    // rom_array[6562] = 32'h00004351;
    // rom_array[6563] = 32'hFFFFFFF1;
    // rom_array[6564] = 32'hFFFFFFF1;
    // rom_array[6565] = 32'h00004359;
    // rom_array[6566] = 32'h00004361;
    // rom_array[6567] = 32'hFFFFFFF1;
    // rom_array[6568] = 32'hFFFFFFF1;
    // rom_array[6569] = 32'h00004369;
    // rom_array[6570] = 32'h00004371;
    // rom_array[6571] = 32'hFFFFFFF1;
    // rom_array[6572] = 32'hFFFFFFF1;
    // rom_array[6573] = 32'h00004379;
    // rom_array[6574] = 32'h00004381;
    // rom_array[6575] = 32'hFFFFFFF1;
    // rom_array[6576] = 32'hFFFFFFF1;
    // rom_array[6577] = 32'h00004389;
    // rom_array[6578] = 32'h00004391;
    // rom_array[6579] = 32'hFFFFFFF1;
    // rom_array[6580] = 32'hFFFFFFF1;
    // rom_array[6581] = 32'h00004399;
    // rom_array[6582] = 32'h000043a1;
    // rom_array[6583] = 32'hFFFFFFF1;
    // rom_array[6584] = 32'hFFFFFFF1;
    // rom_array[6585] = 32'h000043a9;
    // rom_array[6586] = 32'h000043b1;
    // rom_array[6587] = 32'hFFFFFFF0;
    // rom_array[6588] = 32'hFFFFFFF0;
    // rom_array[6589] = 32'h000043b9;
    // rom_array[6590] = 32'h000043c1;
    // rom_array[6591] = 32'hFFFFFFF0;
    // rom_array[6592] = 32'hFFFFFFF0;
    // rom_array[6593] = 32'h000043c9;
    // rom_array[6594] = 32'h000043d1;
    // rom_array[6595] = 32'h000043d9;
    // rom_array[6596] = 32'h000043e1;
    // rom_array[6597] = 32'h000043e9;
    // rom_array[6598] = 32'h000043f1;
    // rom_array[6599] = 32'hFFFFFFF1;
    // rom_array[6600] = 32'hFFFFFFF1;
    // rom_array[6601] = 32'h000043f9;
    // rom_array[6602] = 32'h00004401;
    // rom_array[6603] = 32'h00004409;
    // rom_array[6604] = 32'h00004411;
    // rom_array[6605] = 32'hFFFFFFF1;
    // rom_array[6606] = 32'hFFFFFFF1;
    // rom_array[6607] = 32'hFFFFFFF1;
    // rom_array[6608] = 32'hFFFFFFF1;
    // rom_array[6609] = 32'h00004419;
    // rom_array[6610] = 32'h00004421;
    // rom_array[6611] = 32'h00004429;
    // rom_array[6612] = 32'h00004431;
    // rom_array[6613] = 32'hFFFFFFF1;
    // rom_array[6614] = 32'hFFFFFFF1;
    // rom_array[6615] = 32'hFFFFFFF1;
    // rom_array[6616] = 32'hFFFFFFF1;
    // rom_array[6617] = 32'h00004439;
    // rom_array[6618] = 32'h00004441;
    // rom_array[6619] = 32'h00004449;
    // rom_array[6620] = 32'h00004451;
    // rom_array[6621] = 32'hFFFFFFF1;
    // rom_array[6622] = 32'hFFFFFFF1;
    // rom_array[6623] = 32'hFFFFFFF1;
    // rom_array[6624] = 32'hFFFFFFF1;
    // rom_array[6625] = 32'h00004459;
    // rom_array[6626] = 32'h00004461;
    // rom_array[6627] = 32'hFFFFFFF1;
    // rom_array[6628] = 32'hFFFFFFF1;
    // rom_array[6629] = 32'h00004469;
    // rom_array[6630] = 32'h00004471;
    // rom_array[6631] = 32'hFFFFFFF1;
    // rom_array[6632] = 32'hFFFFFFF1;
    // rom_array[6633] = 32'h00004479;
    // rom_array[6634] = 32'h00004481;
    // rom_array[6635] = 32'h00004489;
    // rom_array[6636] = 32'h00004491;
    // rom_array[6637] = 32'h00004499;
    // rom_array[6638] = 32'h000044a1;
    // rom_array[6639] = 32'hFFFFFFF0;
    // rom_array[6640] = 32'hFFFFFFF0;
    // rom_array[6641] = 32'h000044a9;
    // rom_array[6642] = 32'h000044b1;
    // rom_array[6643] = 32'h000044b9;
    // rom_array[6644] = 32'h000044c1;
    // rom_array[6645] = 32'hFFFFFFF0;
    // rom_array[6646] = 32'hFFFFFFF0;
    // rom_array[6647] = 32'hFFFFFFF0;
    // rom_array[6648] = 32'hFFFFFFF0;
    // rom_array[6649] = 32'h000044c9;
    // rom_array[6650] = 32'h000044d1;
    // rom_array[6651] = 32'h000044d9;
    // rom_array[6652] = 32'h000044e1;
    // rom_array[6653] = 32'hFFFFFFF0;
    // rom_array[6654] = 32'hFFFFFFF0;
    // rom_array[6655] = 32'hFFFFFFF0;
    // rom_array[6656] = 32'hFFFFFFF0;
    // rom_array[6657] = 32'h000044e9;
    // rom_array[6658] = 32'h000044f1;
    // rom_array[6659] = 32'h000044f9;
    // rom_array[6660] = 32'h00004501;
    // rom_array[6661] = 32'hFFFFFFF0;
    // rom_array[6662] = 32'hFFFFFFF0;
    // rom_array[6663] = 32'hFFFFFFF0;
    // rom_array[6664] = 32'hFFFFFFF0;
    // rom_array[6665] = 32'h00004509;
    // rom_array[6666] = 32'h00004511;
    // rom_array[6667] = 32'hFFFFFFF1;
    // rom_array[6668] = 32'hFFFFFFF1;
    // rom_array[6669] = 32'h00004519;
    // rom_array[6670] = 32'h00004521;
    // rom_array[6671] = 32'hFFFFFFF1;
    // rom_array[6672] = 32'hFFFFFFF1;
    // rom_array[6673] = 32'h00004529;
    // rom_array[6674] = 32'h00004531;
    // rom_array[6675] = 32'hFFFFFFF1;
    // rom_array[6676] = 32'hFFFFFFF1;
    // rom_array[6677] = 32'h00004539;
    // rom_array[6678] = 32'h00004541;
    // rom_array[6679] = 32'h00004549;
    // rom_array[6680] = 32'h00004551;
    // rom_array[6681] = 32'hFFFFFFF1;
    // rom_array[6682] = 32'hFFFFFFF1;
    // rom_array[6683] = 32'hFFFFFFF1;
    // rom_array[6684] = 32'hFFFFFFF1;
    // rom_array[6685] = 32'h00004559;
    // rom_array[6686] = 32'h00004561;
    // rom_array[6687] = 32'h00004569;
    // rom_array[6688] = 32'h00004571;
    // rom_array[6689] = 32'h00004579;
    // rom_array[6690] = 32'h00004581;
    // rom_array[6691] = 32'hFFFFFFF0;
    // rom_array[6692] = 32'hFFFFFFF0;
    // rom_array[6693] = 32'h00004589;
    // rom_array[6694] = 32'h00004591;
    // rom_array[6695] = 32'hFFFFFFF0;
    // rom_array[6696] = 32'hFFFFFFF0;
    // rom_array[6697] = 32'h00004599;
    // rom_array[6698] = 32'h000045a1;
    // rom_array[6699] = 32'hFFFFFFF0;
    // rom_array[6700] = 32'hFFFFFFF0;
    // rom_array[6701] = 32'h000045a9;
    // rom_array[6702] = 32'h000045b1;
    // rom_array[6703] = 32'hFFFFFFF0;
    // rom_array[6704] = 32'hFFFFFFF0;
    // rom_array[6705] = 32'h000045b9;
    // rom_array[6706] = 32'h000045c1;
    // rom_array[6707] = 32'h000045c9;
    // rom_array[6708] = 32'h000045d1;
    // rom_array[6709] = 32'h000045d9;
    // rom_array[6710] = 32'h000045e1;
    // rom_array[6711] = 32'hFFFFFFF1;
    // rom_array[6712] = 32'hFFFFFFF1;
    // rom_array[6713] = 32'h000045e9;
    // rom_array[6714] = 32'h000045f1;
    // rom_array[6715] = 32'h000045f9;
    // rom_array[6716] = 32'h00004601;
    // rom_array[6717] = 32'hFFFFFFF1;
    // rom_array[6718] = 32'hFFFFFFF1;
    // rom_array[6719] = 32'hFFFFFFF1;
    // rom_array[6720] = 32'hFFFFFFF1;
    // rom_array[6721] = 32'h00004609;
    // rom_array[6722] = 32'h00004611;
    // rom_array[6723] = 32'h00004619;
    // rom_array[6724] = 32'h00004621;
    // rom_array[6725] = 32'hFFFFFFF1;
    // rom_array[6726] = 32'hFFFFFFF1;
    // rom_array[6727] = 32'hFFFFFFF1;
    // rom_array[6728] = 32'hFFFFFFF1;
    // rom_array[6729] = 32'h00004629;
    // rom_array[6730] = 32'h00004631;
    // rom_array[6731] = 32'h00004639;
    // rom_array[6732] = 32'h00004641;
    // rom_array[6733] = 32'hFFFFFFF1;
    // rom_array[6734] = 32'hFFFFFFF1;
    // rom_array[6735] = 32'h00004649;
    // rom_array[6736] = 32'h00004651;
    // rom_array[6737] = 32'h00004659;
    // rom_array[6738] = 32'h00004661;
    // rom_array[6739] = 32'h00004669;
    // rom_array[6740] = 32'h00004671;
    // rom_array[6741] = 32'h00004679;
    // rom_array[6742] = 32'h00004681;
    // rom_array[6743] = 32'h00004689;
    // rom_array[6744] = 32'h00004691;
    // rom_array[6745] = 32'h00004699;
    // rom_array[6746] = 32'h000046a1;
    // rom_array[6747] = 32'h000046a9;
    // rom_array[6748] = 32'h000046b1;
    // rom_array[6749] = 32'h000046b9;
    // rom_array[6750] = 32'h000046c1;
    // rom_array[6751] = 32'h000046c9;
    // rom_array[6752] = 32'h000046d1;
    // rom_array[6753] = 32'h000046d9;
    // rom_array[6754] = 32'h000046e1;
    // rom_array[6755] = 32'hFFFFFFF1;
    // rom_array[6756] = 32'hFFFFFFF1;
    // rom_array[6757] = 32'h000046e9;
    // rom_array[6758] = 32'h000046f1;
    // rom_array[6759] = 32'hFFFFFFF1;
    // rom_array[6760] = 32'hFFFFFFF1;
    // rom_array[6761] = 32'h000046f9;
    // rom_array[6762] = 32'h00004701;
    // rom_array[6763] = 32'h00004709;
    // rom_array[6764] = 32'h00004711;
    // rom_array[6765] = 32'hFFFFFFF0;
    // rom_array[6766] = 32'hFFFFFFF0;
    // rom_array[6767] = 32'hFFFFFFF0;
    // rom_array[6768] = 32'hFFFFFFF0;
    // rom_array[6769] = 32'h00004719;
    // rom_array[6770] = 32'h00004721;
    // rom_array[6771] = 32'h00004729;
    // rom_array[6772] = 32'h00004731;
    // rom_array[6773] = 32'hFFFFFFF0;
    // rom_array[6774] = 32'hFFFFFFF0;
    // rom_array[6775] = 32'hFFFFFFF0;
    // rom_array[6776] = 32'hFFFFFFF0;
    // rom_array[6777] = 32'hFFFFFFF0;
    // rom_array[6778] = 32'hFFFFFFF0;
    // rom_array[6779] = 32'h00004739;
    // rom_array[6780] = 32'h00004741;
    // rom_array[6781] = 32'hFFFFFFF0;
    // rom_array[6782] = 32'hFFFFFFF0;
    // rom_array[6783] = 32'h00004749;
    // rom_array[6784] = 32'h00004751;
    // rom_array[6785] = 32'h00004759;
    // rom_array[6786] = 32'h00004761;
    // rom_array[6787] = 32'h00004769;
    // rom_array[6788] = 32'h00004771;
    // rom_array[6789] = 32'hFFFFFFF0;
    // rom_array[6790] = 32'hFFFFFFF0;
    // rom_array[6791] = 32'hFFFFFFF0;
    // rom_array[6792] = 32'hFFFFFFF0;
    // rom_array[6793] = 32'h00004779;
    // rom_array[6794] = 32'h00004781;
    // rom_array[6795] = 32'h00004789;
    // rom_array[6796] = 32'h00004791;
    // rom_array[6797] = 32'hFFFFFFF0;
    // rom_array[6798] = 32'hFFFFFFF0;
    // rom_array[6799] = 32'h00004799;
    // rom_array[6800] = 32'h000047a1;
    // rom_array[6801] = 32'h000047a9;
    // rom_array[6802] = 32'h000047b1;
    // rom_array[6803] = 32'h000047b9;
    // rom_array[6804] = 32'h000047c1;
    // rom_array[6805] = 32'hFFFFFFF0;
    // rom_array[6806] = 32'hFFFFFFF0;
    // rom_array[6807] = 32'hFFFFFFF0;
    // rom_array[6808] = 32'hFFFFFFF0;
    // rom_array[6809] = 32'h000047c9;
    // rom_array[6810] = 32'h000047d1;
    // rom_array[6811] = 32'h000047d9;
    // rom_array[6812] = 32'h000047e1;
    // rom_array[6813] = 32'hFFFFFFF0;
    // rom_array[6814] = 32'hFFFFFFF0;
    // rom_array[6815] = 32'hFFFFFFF0;
    // rom_array[6816] = 32'hFFFFFFF0;
    // rom_array[6817] = 32'hFFFFFFF0;
    // rom_array[6818] = 32'hFFFFFFF0;
    // rom_array[6819] = 32'h000047e9;
    // rom_array[6820] = 32'h000047f1;
    // rom_array[6821] = 32'hFFFFFFF0;
    // rom_array[6822] = 32'hFFFFFFF0;
    // rom_array[6823] = 32'h000047f9;
    // rom_array[6824] = 32'h00004801;
    // rom_array[6825] = 32'hFFFFFFF0;
    // rom_array[6826] = 32'hFFFFFFF0;
    // rom_array[6827] = 32'h00004809;
    // rom_array[6828] = 32'h00004811;
    // rom_array[6829] = 32'hFFFFFFF0;
    // rom_array[6830] = 32'hFFFFFFF0;
    // rom_array[6831] = 32'h00004819;
    // rom_array[6832] = 32'h00004821;
    // rom_array[6833] = 32'hFFFFFFF0;
    // rom_array[6834] = 32'hFFFFFFF0;
    // rom_array[6835] = 32'hFFFFFFF0;
    // rom_array[6836] = 32'hFFFFFFF0;
    // rom_array[6837] = 32'hFFFFFFF1;
    // rom_array[6838] = 32'hFFFFFFF1;
    // rom_array[6839] = 32'hFFFFFFF1;
    // rom_array[6840] = 32'hFFFFFFF1;
    // rom_array[6841] = 32'hFFFFFFF0;
    // rom_array[6842] = 32'hFFFFFFF0;
    // rom_array[6843] = 32'hFFFFFFF0;
    // rom_array[6844] = 32'hFFFFFFF0;
    // rom_array[6845] = 32'h00004829;
    // rom_array[6846] = 32'h00004831;
    // rom_array[6847] = 32'hFFFFFFF0;
    // rom_array[6848] = 32'hFFFFFFF0;
    // rom_array[6849] = 32'hFFFFFFF0;
    // rom_array[6850] = 32'hFFFFFFF0;
    // rom_array[6851] = 32'h00004839;
    // rom_array[6852] = 32'h00004841;
    // rom_array[6853] = 32'hFFFFFFF0;
    // rom_array[6854] = 32'hFFFFFFF0;
    // rom_array[6855] = 32'h00004849;
    // rom_array[6856] = 32'h00004851;
    // rom_array[6857] = 32'hFFFFFFF0;
    // rom_array[6858] = 32'hFFFFFFF0;
    // rom_array[6859] = 32'h00004859;
    // rom_array[6860] = 32'h00004861;
    // rom_array[6861] = 32'hFFFFFFF0;
    // rom_array[6862] = 32'hFFFFFFF0;
    // rom_array[6863] = 32'h00004869;
    // rom_array[6864] = 32'h00004871;
    // rom_array[6865] = 32'h00004879;
    // rom_array[6866] = 32'h00004881;
    // rom_array[6867] = 32'h00004889;
    // rom_array[6868] = 32'h00004891;
    // rom_array[6869] = 32'hFFFFFFF1;
    // rom_array[6870] = 32'hFFFFFFF1;
    // rom_array[6871] = 32'hFFFFFFF1;
    // rom_array[6872] = 32'hFFFFFFF1;
    // rom_array[6873] = 32'h00004899;
    // rom_array[6874] = 32'h000048a1;
    // rom_array[6875] = 32'h000048a9;
    // rom_array[6876] = 32'h000048b1;
    // rom_array[6877] = 32'h000048b9;
    // rom_array[6878] = 32'h000048c1;
    // rom_array[6879] = 32'hFFFFFFF1;
    // rom_array[6880] = 32'hFFFFFFF1;
    // rom_array[6881] = 32'h000048c9;
    // rom_array[6882] = 32'h000048d1;
    // rom_array[6883] = 32'h000048d9;
    // rom_array[6884] = 32'h000048e1;
    // rom_array[6885] = 32'hFFFFFFF0;
    // rom_array[6886] = 32'hFFFFFFF0;
    // rom_array[6887] = 32'hFFFFFFF0;
    // rom_array[6888] = 32'hFFFFFFF0;
    // rom_array[6889] = 32'h000048e9;
    // rom_array[6890] = 32'h000048f1;
    // rom_array[6891] = 32'h000048f9;
    // rom_array[6892] = 32'h00004901;
    // rom_array[6893] = 32'h00004909;
    // rom_array[6894] = 32'h00004911;
    // rom_array[6895] = 32'hFFFFFFF0;
    // rom_array[6896] = 32'hFFFFFFF0;
    // rom_array[6897] = 32'hFFFFFFF0;
    // rom_array[6898] = 32'hFFFFFFF0;
    // rom_array[6899] = 32'h00004919;
    // rom_array[6900] = 32'h00004921;
    // rom_array[6901] = 32'hFFFFFFF0;
    // rom_array[6902] = 32'hFFFFFFF0;
    // rom_array[6903] = 32'h00004929;
    // rom_array[6904] = 32'h00004931;
    // rom_array[6905] = 32'hFFFFFFF0;
    // rom_array[6906] = 32'hFFFFFFF0;
    // rom_array[6907] = 32'h00004939;
    // rom_array[6908] = 32'h00004941;
    // rom_array[6909] = 32'hFFFFFFF0;
    // rom_array[6910] = 32'hFFFFFFF0;
    // rom_array[6911] = 32'h00004949;
    // rom_array[6912] = 32'h00004951;
    // rom_array[6913] = 32'h00004959;
    // rom_array[6914] = 32'h00004961;
    // rom_array[6915] = 32'h00004969;
    // rom_array[6916] = 32'h00004971;
    // rom_array[6917] = 32'h00004979;
    // rom_array[6918] = 32'h00004981;
    // rom_array[6919] = 32'hFFFFFFF1;
    // rom_array[6920] = 32'hFFFFFFF1;
    // rom_array[6921] = 32'h00004989;
    // rom_array[6922] = 32'h00004991;
    // rom_array[6923] = 32'h00004999;
    // rom_array[6924] = 32'h000049a1;
    // rom_array[6925] = 32'hFFFFFFF1;
    // rom_array[6926] = 32'hFFFFFFF1;
    // rom_array[6927] = 32'hFFFFFFF1;
    // rom_array[6928] = 32'hFFFFFFF1;
    // rom_array[6929] = 32'h000049a9;
    // rom_array[6930] = 32'h000049b1;
    // rom_array[6931] = 32'hFFFFFFF1;
    // rom_array[6932] = 32'hFFFFFFF1;
    // rom_array[6933] = 32'h000049b9;
    // rom_array[6934] = 32'h000049c1;
    // rom_array[6935] = 32'hFFFFFFF1;
    // rom_array[6936] = 32'hFFFFFFF1;
    // rom_array[6937] = 32'h000049c9;
    // rom_array[6938] = 32'h000049d1;
    // rom_array[6939] = 32'h000049d9;
    // rom_array[6940] = 32'h000049e1;
    // rom_array[6941] = 32'hFFFFFFF0;
    // rom_array[6942] = 32'hFFFFFFF0;
    // rom_array[6943] = 32'hFFFFFFF0;
    // rom_array[6944] = 32'hFFFFFFF0;
    // rom_array[6945] = 32'h000049e9;
    // rom_array[6946] = 32'h000049f1;
    // rom_array[6947] = 32'h000049f9;
    // rom_array[6948] = 32'h00004a01;
    // rom_array[6949] = 32'hFFFFFFF0;
    // rom_array[6950] = 32'hFFFFFFF0;
    // rom_array[6951] = 32'hFFFFFFF0;
    // rom_array[6952] = 32'hFFFFFFF0;
    // rom_array[6953] = 32'h00004a09;
    // rom_array[6954] = 32'h00004a11;
    // rom_array[6955] = 32'h00004a19;
    // rom_array[6956] = 32'h00004a21;
    // rom_array[6957] = 32'hFFFFFFF1;
    // rom_array[6958] = 32'hFFFFFFF1;
    // rom_array[6959] = 32'hFFFFFFF1;
    // rom_array[6960] = 32'hFFFFFFF1;
    // rom_array[6961] = 32'h00004a29;
    // rom_array[6962] = 32'h00004a31;
    // rom_array[6963] = 32'h00004a39;
    // rom_array[6964] = 32'h00004a41;
    // rom_array[6965] = 32'hFFFFFFF1;
    // rom_array[6966] = 32'hFFFFFFF1;
    // rom_array[6967] = 32'h00004a49;
    // rom_array[6968] = 32'h00004a51;
    // rom_array[6969] = 32'hFFFFFFF0;
    // rom_array[6970] = 32'hFFFFFFF0;
    // rom_array[6971] = 32'h00004a59;
    // rom_array[6972] = 32'h00004a61;
    // rom_array[6973] = 32'hFFFFFFF0;
    // rom_array[6974] = 32'hFFFFFFF0;
    // rom_array[6975] = 32'h00004a69;
    // rom_array[6976] = 32'h00004a71;
    // rom_array[6977] = 32'h00004a79;
    // rom_array[6978] = 32'h00004a81;
    // rom_array[6979] = 32'h00004a89;
    // rom_array[6980] = 32'h00004a91;
    // rom_array[6981] = 32'hFFFFFFF1;
    // rom_array[6982] = 32'hFFFFFFF1;
    // rom_array[6983] = 32'hFFFFFFF1;
    // rom_array[6984] = 32'hFFFFFFF1;
    // rom_array[6985] = 32'h00004a99;
    // rom_array[6986] = 32'h00004aa1;
    // rom_array[6987] = 32'h00004aa9;
    // rom_array[6988] = 32'h00004ab1;
    // rom_array[6989] = 32'hFFFFFFF1;
    // rom_array[6990] = 32'hFFFFFFF1;
    // rom_array[6991] = 32'hFFFFFFF1;
    // rom_array[6992] = 32'hFFFFFFF1;
    // rom_array[6993] = 32'hFFFFFFF1;
    // rom_array[6994] = 32'hFFFFFFF1;
    // rom_array[6995] = 32'hFFFFFFF1;
    // rom_array[6996] = 32'hFFFFFFF1;
    // rom_array[6997] = 32'h00004ab9;
    // rom_array[6998] = 32'h00004ac1;
    // rom_array[6999] = 32'h00004ac9;
    // rom_array[7000] = 32'h00004ad1;
    // rom_array[7001] = 32'hFFFFFFF1;
    // rom_array[7002] = 32'hFFFFFFF1;
    // rom_array[7003] = 32'hFFFFFFF1;
    // rom_array[7004] = 32'hFFFFFFF1;
    // rom_array[7005] = 32'h00004ad9;
    // rom_array[7006] = 32'h00004ae1;
    // rom_array[7007] = 32'h00004ae9;
    // rom_array[7008] = 32'h00004af1;
    // rom_array[7009] = 32'h00004af9;
    // rom_array[7010] = 32'h00004b01;
    // rom_array[7011] = 32'h00004b09;
    // rom_array[7012] = 32'h00004b11;
    // rom_array[7013] = 32'hFFFFFFF0;
    // rom_array[7014] = 32'hFFFFFFF0;
    // rom_array[7015] = 32'hFFFFFFF0;
    // rom_array[7016] = 32'hFFFFFFF0;
    // rom_array[7017] = 32'h00004b19;
    // rom_array[7018] = 32'h00004b21;
    // rom_array[7019] = 32'h00004b29;
    // rom_array[7020] = 32'h00004b31;
    // rom_array[7021] = 32'hFFFFFFF0;
    // rom_array[7022] = 32'hFFFFFFF0;
    // rom_array[7023] = 32'hFFFFFFF0;
    // rom_array[7024] = 32'hFFFFFFF0;
    // rom_array[7025] = 32'h00004b39;
    // rom_array[7026] = 32'h00004b41;
    // rom_array[7027] = 32'h00004b49;
    // rom_array[7028] = 32'h00004b51;
    // rom_array[7029] = 32'hFFFFFFF0;
    // rom_array[7030] = 32'hFFFFFFF0;
    // rom_array[7031] = 32'hFFFFFFF0;
    // rom_array[7032] = 32'hFFFFFFF0;
    // rom_array[7033] = 32'h00004b59;
    // rom_array[7034] = 32'h00004b61;
    // rom_array[7035] = 32'h00004b69;
    // rom_array[7036] = 32'h00004b71;
    // rom_array[7037] = 32'hFFFFFFF0;
    // rom_array[7038] = 32'hFFFFFFF0;
    // rom_array[7039] = 32'hFFFFFFF0;
    // rom_array[7040] = 32'hFFFFFFF0;
    // rom_array[7041] = 32'h00004b79;
    // rom_array[7042] = 32'h00004b81;
    // rom_array[7043] = 32'h00004b89;
    // rom_array[7044] = 32'h00004b91;
    // rom_array[7045] = 32'h00004b99;
    // rom_array[7046] = 32'h00004ba1;
    // rom_array[7047] = 32'hFFFFFFF1;
    // rom_array[7048] = 32'hFFFFFFF1;
    // rom_array[7049] = 32'h00004ba9;
    // rom_array[7050] = 32'h00004bb1;
    // rom_array[7051] = 32'h00004bb9;
    // rom_array[7052] = 32'h00004bc1;
    // rom_array[7053] = 32'hFFFFFFF1;
    // rom_array[7054] = 32'hFFFFFFF1;
    // rom_array[7055] = 32'hFFFFFFF1;
    // rom_array[7056] = 32'hFFFFFFF1;
    // rom_array[7057] = 32'h00004bc9;
    // rom_array[7058] = 32'h00004bd1;
    // rom_array[7059] = 32'hFFFFFFF1;
    // rom_array[7060] = 32'hFFFFFFF1;
    // rom_array[7061] = 32'h00004bd9;
    // rom_array[7062] = 32'h00004be1;
    // rom_array[7063] = 32'hFFFFFFF1;
    // rom_array[7064] = 32'hFFFFFFF1;
    // rom_array[7065] = 32'h00004be9;
    // rom_array[7066] = 32'h00004bf1;
    // rom_array[7067] = 32'h00004bf9;
    // rom_array[7068] = 32'h00004c01;
    // rom_array[7069] = 32'hFFFFFFF0;
    // rom_array[7070] = 32'hFFFFFFF0;
    // rom_array[7071] = 32'hFFFFFFF0;
    // rom_array[7072] = 32'hFFFFFFF0;
    // rom_array[7073] = 32'h00004c09;
    // rom_array[7074] = 32'h00004c11;
    // rom_array[7075] = 32'h00004c19;
    // rom_array[7076] = 32'h00004c21;
    // rom_array[7077] = 32'hFFFFFFF0;
    // rom_array[7078] = 32'hFFFFFFF0;
    // rom_array[7079] = 32'hFFFFFFF0;
    // rom_array[7080] = 32'hFFFFFFF0;
    // rom_array[7081] = 32'h00004c29;
    // rom_array[7082] = 32'h00004c31;
    // rom_array[7083] = 32'h00004c39;
    // rom_array[7084] = 32'h00004c41;
    // rom_array[7085] = 32'hFFFFFFF1;
    // rom_array[7086] = 32'hFFFFFFF1;
    // rom_array[7087] = 32'hFFFFFFF1;
    // rom_array[7088] = 32'hFFFFFFF1;
    // rom_array[7089] = 32'h00004c49;
    // rom_array[7090] = 32'h00004c51;
    // rom_array[7091] = 32'h00004c59;
    // rom_array[7092] = 32'h00004c61;
    // rom_array[7093] = 32'hFFFFFFF1;
    // rom_array[7094] = 32'hFFFFFFF1;
    // rom_array[7095] = 32'hFFFFFFF1;
    // rom_array[7096] = 32'hFFFFFFF1;
    // rom_array[7097] = 32'h00004c69;
    // rom_array[7098] = 32'h00004c71;
    // rom_array[7099] = 32'h00004c79;
    // rom_array[7100] = 32'h00004c81;
    // rom_array[7101] = 32'hFFFFFFF1;
    // rom_array[7102] = 32'hFFFFFFF1;
    // rom_array[7103] = 32'hFFFFFFF1;
    // rom_array[7104] = 32'hFFFFFFF1;
    // rom_array[7105] = 32'h00004c89;
    // rom_array[7106] = 32'h00004c91;
    // rom_array[7107] = 32'h00004c99;
    // rom_array[7108] = 32'h00004ca1;
    // rom_array[7109] = 32'hFFFFFFF1;
    // rom_array[7110] = 32'hFFFFFFF1;
    // rom_array[7111] = 32'hFFFFFFF1;
    // rom_array[7112] = 32'hFFFFFFF1;
    // rom_array[7113] = 32'h00004ca9;
    // rom_array[7114] = 32'h00004cb1;
    // rom_array[7115] = 32'h00004cb9;
    // rom_array[7116] = 32'h00004cc1;
    // rom_array[7117] = 32'hFFFFFFF0;
    // rom_array[7118] = 32'hFFFFFFF0;
    // rom_array[7119] = 32'hFFFFFFF0;
    // rom_array[7120] = 32'hFFFFFFF0;
    // rom_array[7121] = 32'h00004cc9;
    // rom_array[7122] = 32'h00004cd1;
    // rom_array[7123] = 32'h00004cd9;
    // rom_array[7124] = 32'h00004ce1;
    // rom_array[7125] = 32'hFFFFFFF0;
    // rom_array[7126] = 32'hFFFFFFF0;
    // rom_array[7127] = 32'hFFFFFFF0;
    // rom_array[7128] = 32'hFFFFFFF0;
    // rom_array[7129] = 32'h00004ce9;
    // rom_array[7130] = 32'h00004cf1;
    // rom_array[7131] = 32'h00004cf9;
    // rom_array[7132] = 32'h00004d01;
    // rom_array[7133] = 32'h00004d09;
    // rom_array[7134] = 32'h00004d11;
    // rom_array[7135] = 32'hFFFFFFF1;
    // rom_array[7136] = 32'hFFFFFFF1;
    // rom_array[7137] = 32'h00004d19;
    // rom_array[7138] = 32'h00004d21;
    // rom_array[7139] = 32'h00004d29;
    // rom_array[7140] = 32'h00004d31;
    // rom_array[7141] = 32'hFFFFFFF1;
    // rom_array[7142] = 32'hFFFFFFF1;
    // rom_array[7143] = 32'hFFFFFFF1;
    // rom_array[7144] = 32'hFFFFFFF1;
    // rom_array[7145] = 32'h00004d39;
    // rom_array[7146] = 32'h00004d41;
    // rom_array[7147] = 32'hFFFFFFF1;
    // rom_array[7148] = 32'hFFFFFFF1;
    // rom_array[7149] = 32'h00004d49;
    // rom_array[7150] = 32'h00004d51;
    // rom_array[7151] = 32'hFFFFFFF1;
    // rom_array[7152] = 32'hFFFFFFF1;
    // rom_array[7153] = 32'h00004d59;
    // rom_array[7154] = 32'h00004d61;
    // rom_array[7155] = 32'hFFFFFFF1;
    // rom_array[7156] = 32'hFFFFFFF1;
    // rom_array[7157] = 32'h00004d69;
    // rom_array[7158] = 32'h00004d71;
    // rom_array[7159] = 32'hFFFFFFF1;
    // rom_array[7160] = 32'hFFFFFFF1;
    // rom_array[7161] = 32'h00004d79;
    // rom_array[7162] = 32'h00004d81;
    // rom_array[7163] = 32'hFFFFFFF1;
    // rom_array[7164] = 32'hFFFFFFF1;
    // rom_array[7165] = 32'h00004d89;
    // rom_array[7166] = 32'h00004d91;
    // rom_array[7167] = 32'hFFFFFFF1;
    // rom_array[7168] = 32'hFFFFFFF1;
    // rom_array[7169] = 32'hFFFFFFF0;
    // rom_array[7170] = 32'hFFFFFFF0;
    // rom_array[7171] = 32'hFFFFFFF0;
    // rom_array[7172] = 32'hFFFFFFF0;
    // rom_array[7173] = 32'hFFFFFFF0;
    // rom_array[7174] = 32'hFFFFFFF0;
    // rom_array[7175] = 32'h00004d99;
    // rom_array[7176] = 32'h00004da1;
    // rom_array[7177] = 32'h00004da9;
    // rom_array[7178] = 32'h00004db1;
    // rom_array[7179] = 32'h00004db9;
    // rom_array[7180] = 32'h00004dc1;
    // rom_array[7181] = 32'hFFFFFFF0;
    // rom_array[7182] = 32'hFFFFFFF0;
    // rom_array[7183] = 32'hFFFFFFF0;
    // rom_array[7184] = 32'hFFFFFFF0;
    // rom_array[7185] = 32'h00004dc9;
    // rom_array[7186] = 32'h00004dd1;
    // rom_array[7187] = 32'h00004dd9;
    // rom_array[7188] = 32'h00004de1;
    // rom_array[7189] = 32'hFFFFFFF0;
    // rom_array[7190] = 32'hFFFFFFF0;
    // rom_array[7191] = 32'h00004de9;
    // rom_array[7192] = 32'h00004df1;
    // rom_array[7193] = 32'hFFFFFFF0;
    // rom_array[7194] = 32'hFFFFFFF0;
    // rom_array[7195] = 32'h00004df9;
    // rom_array[7196] = 32'h00004e01;
    // rom_array[7197] = 32'hFFFFFFF0;
    // rom_array[7198] = 32'hFFFFFFF0;
    // rom_array[7199] = 32'h00004e09;
    // rom_array[7200] = 32'h00004e11;
    // rom_array[7201] = 32'h00004e19;
    // rom_array[7202] = 32'h00004e21;
    // rom_array[7203] = 32'h00004e29;
    // rom_array[7204] = 32'h00004e31;
    // rom_array[7205] = 32'h00004e39;
    // rom_array[7206] = 32'h00004e41;
    // rom_array[7207] = 32'hFFFFFFF1;
    // rom_array[7208] = 32'hFFFFFFF1;
    // rom_array[7209] = 32'h00004e49;
    // rom_array[7210] = 32'h00004e51;
    // rom_array[7211] = 32'h00004e59;
    // rom_array[7212] = 32'h00004e61;
    // rom_array[7213] = 32'hFFFFFFF1;
    // rom_array[7214] = 32'hFFFFFFF1;
    // rom_array[7215] = 32'hFFFFFFF1;
    // rom_array[7216] = 32'hFFFFFFF1;
    // rom_array[7217] = 32'h00004e69;
    // rom_array[7218] = 32'h00004e71;
    // rom_array[7219] = 32'hFFFFFFF1;
    // rom_array[7220] = 32'hFFFFFFF1;
    // rom_array[7221] = 32'h00004e79;
    // rom_array[7222] = 32'h00004e81;
    // rom_array[7223] = 32'hFFFFFFF1;
    // rom_array[7224] = 32'hFFFFFFF1;
    // rom_array[7225] = 32'h00004e89;
    // rom_array[7226] = 32'h00004e91;
    // rom_array[7227] = 32'h00004e99;
    // rom_array[7228] = 32'h00004ea1;
    // rom_array[7229] = 32'h00004ea9;
    // rom_array[7230] = 32'h00004eb1;
    // rom_array[7231] = 32'hFFFFFFF1;
    // rom_array[7232] = 32'hFFFFFFF1;
    // rom_array[7233] = 32'h00004eb9;
    // rom_array[7234] = 32'h00004ec1;
    // rom_array[7235] = 32'h00004ec9;
    // rom_array[7236] = 32'h00004ed1;
    // rom_array[7237] = 32'hFFFFFFF1;
    // rom_array[7238] = 32'hFFFFFFF1;
    // rom_array[7239] = 32'hFFFFFFF1;
    // rom_array[7240] = 32'hFFFFFFF1;
    // rom_array[7241] = 32'h00004ed9;
    // rom_array[7242] = 32'h00004ee1;
    // rom_array[7243] = 32'h00004ee9;
    // rom_array[7244] = 32'h00004ef1;
    // rom_array[7245] = 32'hFFFFFFF1;
    // rom_array[7246] = 32'hFFFFFFF1;
    // rom_array[7247] = 32'hFFFFFFF1;
    // rom_array[7248] = 32'hFFFFFFF1;
    // rom_array[7249] = 32'h00004ef9;
    // rom_array[7250] = 32'h00004f01;
    // rom_array[7251] = 32'h00004f09;
    // rom_array[7252] = 32'h00004f11;
    // rom_array[7253] = 32'hFFFFFFF1;
    // rom_array[7254] = 32'hFFFFFFF1;
    // rom_array[7255] = 32'hFFFFFFF1;
    // rom_array[7256] = 32'hFFFFFFF1;
    // rom_array[7257] = 32'h00004f19;
    // rom_array[7258] = 32'h00004f21;
    // rom_array[7259] = 32'h00004f29;
    // rom_array[7260] = 32'h00004f31;
    // rom_array[7261] = 32'hFFFFFFF1;
    // rom_array[7262] = 32'hFFFFFFF1;
    // rom_array[7263] = 32'hFFFFFFF1;
    // rom_array[7264] = 32'hFFFFFFF1;
    // rom_array[7265] = 32'h00004f39;
    // rom_array[7266] = 32'h00004f41;
    // rom_array[7267] = 32'h00004f49;
    // rom_array[7268] = 32'h00004f51;
    // rom_array[7269] = 32'hFFFFFFF1;
    // rom_array[7270] = 32'hFFFFFFF1;
    // rom_array[7271] = 32'hFFFFFFF1;
    // rom_array[7272] = 32'hFFFFFFF1;
    // rom_array[7273] = 32'h00004f59;
    // rom_array[7274] = 32'h00004f61;
    // rom_array[7275] = 32'h00004f69;
    // rom_array[7276] = 32'h00004f71;
    // rom_array[7277] = 32'h00004f79;
    // rom_array[7278] = 32'h00004f81;
    // rom_array[7279] = 32'hFFFFFFF0;
    // rom_array[7280] = 32'hFFFFFFF0;
    // rom_array[7281] = 32'h00004f89;
    // rom_array[7282] = 32'h00004f91;
    // rom_array[7283] = 32'h00004f99;
    // rom_array[7284] = 32'h00004fa1;
    // rom_array[7285] = 32'hFFFFFFF0;
    // rom_array[7286] = 32'hFFFFFFF0;
    // rom_array[7287] = 32'hFFFFFFF0;
    // rom_array[7288] = 32'hFFFFFFF0;
    // rom_array[7289] = 32'h00004fa9;
    // rom_array[7290] = 32'h00004fb1;
    // rom_array[7291] = 32'h00004fb9;
    // rom_array[7292] = 32'h00004fc1;
    // rom_array[7293] = 32'hFFFFFFF0;
    // rom_array[7294] = 32'hFFFFFFF0;
    // rom_array[7295] = 32'h00004fc9;
    // rom_array[7296] = 32'h00004fd1;
    // rom_array[7297] = 32'h00004fd9;
    // rom_array[7298] = 32'h00004fe1;
    // rom_array[7299] = 32'h00004fe9;
    // rom_array[7300] = 32'h00004ff1;
    // rom_array[7301] = 32'hFFFFFFF1;
    // rom_array[7302] = 32'hFFFFFFF1;
    // rom_array[7303] = 32'hFFFFFFF1;
    // rom_array[7304] = 32'hFFFFFFF1;
    // rom_array[7305] = 32'h00004ff9;
    // rom_array[7306] = 32'h00005001;
    // rom_array[7307] = 32'hFFFFFFF1;
    // rom_array[7308] = 32'hFFFFFFF1;
    // rom_array[7309] = 32'h00005009;
    // rom_array[7310] = 32'h00005011;
    // rom_array[7311] = 32'hFFFFFFF1;
    // rom_array[7312] = 32'hFFFFFFF1;
    // rom_array[7313] = 32'h00005019;
    // rom_array[7314] = 32'h00005021;
    // rom_array[7315] = 32'hFFFFFFF1;
    // rom_array[7316] = 32'hFFFFFFF1;
    // rom_array[7317] = 32'h00005029;
    // rom_array[7318] = 32'h00005031;
    // rom_array[7319] = 32'hFFFFFFF1;
    // rom_array[7320] = 32'hFFFFFFF1;
    // rom_array[7321] = 32'h00005039;
    // rom_array[7322] = 32'h00005041;
    // rom_array[7323] = 32'hFFFFFFF1;
    // rom_array[7324] = 32'hFFFFFFF1;
    // rom_array[7325] = 32'h00005049;
    // rom_array[7326] = 32'h00005051;
    // rom_array[7327] = 32'hFFFFFFF1;
    // rom_array[7328] = 32'hFFFFFFF1;
    // rom_array[7329] = 32'h00005059;
    // rom_array[7330] = 32'h00005061;
    // rom_array[7331] = 32'hFFFFFFF1;
    // rom_array[7332] = 32'hFFFFFFF1;
    // rom_array[7333] = 32'h00005069;
    // rom_array[7334] = 32'h00005071;
    // rom_array[7335] = 32'hFFFFFFF1;
    // rom_array[7336] = 32'hFFFFFFF1;
    // rom_array[7337] = 32'h00005079;
    // rom_array[7338] = 32'h00005081;
    // rom_array[7339] = 32'hFFFFFFF0;
    // rom_array[7340] = 32'hFFFFFFF0;
    // rom_array[7341] = 32'h00005089;
    // rom_array[7342] = 32'h00005091;
    // rom_array[7343] = 32'hFFFFFFF0;
    // rom_array[7344] = 32'hFFFFFFF0;
    // rom_array[7345] = 32'h00005099;
    // rom_array[7346] = 32'h000050a1;
    // rom_array[7347] = 32'hFFFFFFF0;
    // rom_array[7348] = 32'hFFFFFFF0;
    // rom_array[7349] = 32'h000050a9;
    // rom_array[7350] = 32'h000050b1;
    // rom_array[7351] = 32'hFFFFFFF0;
    // rom_array[7352] = 32'hFFFFFFF0;
    // rom_array[7353] = 32'hFFFFFFF0;
    // rom_array[7354] = 32'hFFFFFFF0;
    // rom_array[7355] = 32'h000050b9;
    // rom_array[7356] = 32'h000050c1;
    // rom_array[7357] = 32'hFFFFFFF0;
    // rom_array[7358] = 32'hFFFFFFF0;
    // rom_array[7359] = 32'h000050c9;
    // rom_array[7360] = 32'h000050d1;
    // rom_array[7361] = 32'hFFFFFFF0;
    // rom_array[7362] = 32'hFFFFFFF0;
    // rom_array[7363] = 32'h000050d9;
    // rom_array[7364] = 32'h000050e1;
    // rom_array[7365] = 32'hFFFFFFF0;
    // rom_array[7366] = 32'hFFFFFFF0;
    // rom_array[7367] = 32'h000050e9;
    // rom_array[7368] = 32'h000050f1;
    // rom_array[7369] = 32'h000050f9;
    // rom_array[7370] = 32'h00005101;
    // rom_array[7371] = 32'hFFFFFFF0;
    // rom_array[7372] = 32'hFFFFFFF0;
    // rom_array[7373] = 32'h00005109;
    // rom_array[7374] = 32'h00005111;
    // rom_array[7375] = 32'hFFFFFFF0;
    // rom_array[7376] = 32'hFFFFFFF0;
    // rom_array[7377] = 32'h00005119;
    // rom_array[7378] = 32'h00005121;
    // rom_array[7379] = 32'hFFFFFFF0;
    // rom_array[7380] = 32'hFFFFFFF0;
    // rom_array[7381] = 32'h00005129;
    // rom_array[7382] = 32'h00005131;
    // rom_array[7383] = 32'hFFFFFFF0;
    // rom_array[7384] = 32'hFFFFFFF0;
    // rom_array[7385] = 32'hFFFFFFF0;
    // rom_array[7386] = 32'hFFFFFFF0;
    // rom_array[7387] = 32'h00005139;
    // rom_array[7388] = 32'h00005141;
    // rom_array[7389] = 32'hFFFFFFF0;
    // rom_array[7390] = 32'hFFFFFFF0;
    // rom_array[7391] = 32'h00005149;
    // rom_array[7392] = 32'h00005151;
    // rom_array[7393] = 32'hFFFFFFF0;
    // rom_array[7394] = 32'hFFFFFFF0;
    // rom_array[7395] = 32'h00005159;
    // rom_array[7396] = 32'h00005161;
    // rom_array[7397] = 32'hFFFFFFF0;
    // rom_array[7398] = 32'hFFFFFFF0;
    // rom_array[7399] = 32'h00005169;
    // rom_array[7400] = 32'h00005171;
    // rom_array[7401] = 32'hFFFFFFF0;
    // rom_array[7402] = 32'hFFFFFFF0;
    // rom_array[7403] = 32'hFFFFFFF0;
    // rom_array[7404] = 32'hFFFFFFF0;
    // rom_array[7405] = 32'h00005179;
    // rom_array[7406] = 32'h00005181;
    // rom_array[7407] = 32'h00005189;
    // rom_array[7408] = 32'h00005191;
    // rom_array[7409] = 32'h00005199;
    // rom_array[7410] = 32'h000051a1;
    // rom_array[7411] = 32'hFFFFFFF1;
    // rom_array[7412] = 32'hFFFFFFF1;
    // rom_array[7413] = 32'h000051a9;
    // rom_array[7414] = 32'h000051b1;
    // rom_array[7415] = 32'hFFFFFFF1;
    // rom_array[7416] = 32'hFFFFFFF1;
    // rom_array[7417] = 32'hFFFFFFF0;
    // rom_array[7418] = 32'hFFFFFFF0;
    // rom_array[7419] = 32'hFFFFFFF0;
    // rom_array[7420] = 32'hFFFFFFF0;
    // rom_array[7421] = 32'h000051b9;
    // rom_array[7422] = 32'h000051c1;
    // rom_array[7423] = 32'h000051c9;
    // rom_array[7424] = 32'h000051d1;
    // rom_array[7425] = 32'hFFFFFFF0;
    // rom_array[7426] = 32'hFFFFFFF0;
    // rom_array[7427] = 32'hFFFFFFF0;
    // rom_array[7428] = 32'hFFFFFFF0;
    // rom_array[7429] = 32'h000051d9;
    // rom_array[7430] = 32'h000051e1;
    // rom_array[7431] = 32'hFFFFFFF0;
    // rom_array[7432] = 32'hFFFFFFF0;
    // rom_array[7433] = 32'h000051e9;
    // rom_array[7434] = 32'h000051f1;
    // rom_array[7435] = 32'hFFFFFFF0;
    // rom_array[7436] = 32'hFFFFFFF0;
    // rom_array[7437] = 32'h000051f9;
    // rom_array[7438] = 32'h00005201;
    // rom_array[7439] = 32'hFFFFFFF0;
    // rom_array[7440] = 32'hFFFFFFF0;
    // rom_array[7441] = 32'h00005209;
    // rom_array[7442] = 32'h00005211;
    // rom_array[7443] = 32'h00005219;
    // rom_array[7444] = 32'h00005221;
    // rom_array[7445] = 32'hFFFFFFF1;
    // rom_array[7446] = 32'hFFFFFFF1;
    // rom_array[7447] = 32'hFFFFFFF1;
    // rom_array[7448] = 32'hFFFFFFF1;
    // rom_array[7449] = 32'h00005229;
    // rom_array[7450] = 32'h00005231;
    // rom_array[7451] = 32'h00005239;
    // rom_array[7452] = 32'h00005241;
    // rom_array[7453] = 32'hFFFFFFF1;
    // rom_array[7454] = 32'hFFFFFFF1;
    // rom_array[7455] = 32'hFFFFFFF1;
    // rom_array[7456] = 32'hFFFFFFF1;
    // rom_array[7457] = 32'h00005249;
    // rom_array[7458] = 32'h00005251;
    // rom_array[7459] = 32'hFFFFFFF1;
    // rom_array[7460] = 32'hFFFFFFF1;
    // rom_array[7461] = 32'h00005259;
    // rom_array[7462] = 32'h00005261;
    // rom_array[7463] = 32'hFFFFFFF1;
    // rom_array[7464] = 32'hFFFFFFF1;
    // rom_array[7465] = 32'h00005269;
    // rom_array[7466] = 32'h00005271;
    // rom_array[7467] = 32'h00005279;
    // rom_array[7468] = 32'h00005281;
    // rom_array[7469] = 32'hFFFFFFF1;
    // rom_array[7470] = 32'hFFFFFFF1;
    // rom_array[7471] = 32'hFFFFFFF1;
    // rom_array[7472] = 32'hFFFFFFF1;
    // rom_array[7473] = 32'h00005289;
    // rom_array[7474] = 32'h00005291;
    // rom_array[7475] = 32'hFFFFFFF1;
    // rom_array[7476] = 32'hFFFFFFF1;
    // rom_array[7477] = 32'h00005299;
    // rom_array[7478] = 32'h000052a1;
    // rom_array[7479] = 32'hFFFFFFF1;
    // rom_array[7480] = 32'hFFFFFFF1;
    // rom_array[7481] = 32'h000052a9;
    // rom_array[7482] = 32'h000052b1;
    // rom_array[7483] = 32'h000052b9;
    // rom_array[7484] = 32'h000052c1;
    // rom_array[7485] = 32'hFFFFFFF0;
    // rom_array[7486] = 32'hFFFFFFF0;
    // rom_array[7487] = 32'hFFFFFFF0;
    // rom_array[7488] = 32'hFFFFFFF0;
    // rom_array[7489] = 32'h000052c9;
    // rom_array[7490] = 32'h000052d1;
    // rom_array[7491] = 32'h000052d9;
    // rom_array[7492] = 32'h000052e1;
    // rom_array[7493] = 32'hFFFFFFF0;
    // rom_array[7494] = 32'hFFFFFFF0;
    // rom_array[7495] = 32'hFFFFFFF0;
    // rom_array[7496] = 32'hFFFFFFF0;
    // rom_array[7497] = 32'h000052e9;
    // rom_array[7498] = 32'h000052f1;
    // rom_array[7499] = 32'hFFFFFFF1;
    // rom_array[7500] = 32'hFFFFFFF1;
    // rom_array[7501] = 32'h000052f9;
    // rom_array[7502] = 32'h00005301;
    // rom_array[7503] = 32'hFFFFFFF1;
    // rom_array[7504] = 32'hFFFFFFF1;
    // rom_array[7505] = 32'h00005309;
    // rom_array[7506] = 32'h00005311;
    // rom_array[7507] = 32'h00005319;
    // rom_array[7508] = 32'h00005321;
    // rom_array[7509] = 32'hFFFFFFF0;
    // rom_array[7510] = 32'hFFFFFFF0;
    // rom_array[7511] = 32'hFFFFFFF0;
    // rom_array[7512] = 32'hFFFFFFF0;
    // rom_array[7513] = 32'h00005329;
    // rom_array[7514] = 32'h00005331;
    // rom_array[7515] = 32'hFFFFFFF1;
    // rom_array[7516] = 32'hFFFFFFF1;
    // rom_array[7517] = 32'h00005339;
    // rom_array[7518] = 32'h00005341;
    // rom_array[7519] = 32'hFFFFFFF1;
    // rom_array[7520] = 32'hFFFFFFF1;
    // rom_array[7521] = 32'h00005349;
    // rom_array[7522] = 32'h00005351;
    // rom_array[7523] = 32'hFFFFFFF0;
    // rom_array[7524] = 32'hFFFFFFF0;
    // rom_array[7525] = 32'h00005359;
    // rom_array[7526] = 32'h00005361;
    // rom_array[7527] = 32'hFFFFFFF0;
    // rom_array[7528] = 32'hFFFFFFF0;
    // rom_array[7529] = 32'h00005369;
    // rom_array[7530] = 32'h00005371;
    // rom_array[7531] = 32'hFFFFFFF0;
    // rom_array[7532] = 32'hFFFFFFF0;
    // rom_array[7533] = 32'h00005379;
    // rom_array[7534] = 32'h00005381;
    // rom_array[7535] = 32'hFFFFFFF0;
    // rom_array[7536] = 32'hFFFFFFF0;
    // rom_array[7537] = 32'h00005389;
    // rom_array[7538] = 32'h00005391;
    // rom_array[7539] = 32'hFFFFFFF0;
    // rom_array[7540] = 32'hFFFFFFF0;
    // rom_array[7541] = 32'h00005399;
    // rom_array[7542] = 32'h000053a1;
    // rom_array[7543] = 32'hFFFFFFF0;
    // rom_array[7544] = 32'hFFFFFFF0;
    // rom_array[7545] = 32'h000053a9;
    // rom_array[7546] = 32'h000053b1;
    // rom_array[7547] = 32'hFFFFFFF0;
    // rom_array[7548] = 32'hFFFFFFF0;
    // rom_array[7549] = 32'h000053b9;
    // rom_array[7550] = 32'h000053c1;
    // rom_array[7551] = 32'hFFFFFFF0;
    // rom_array[7552] = 32'hFFFFFFF0;
    // rom_array[7553] = 32'h000053c9;
    // rom_array[7554] = 32'h000053d1;
    // rom_array[7555] = 32'hFFFFFFF1;
    // rom_array[7556] = 32'hFFFFFFF1;
    // rom_array[7557] = 32'h000053d9;
    // rom_array[7558] = 32'h000053e1;
    // rom_array[7559] = 32'hFFFFFFF1;
    // rom_array[7560] = 32'hFFFFFFF1;
    // rom_array[7561] = 32'h000053e9;
    // rom_array[7562] = 32'h000053f1;
    // rom_array[7563] = 32'hFFFFFFF1;
    // rom_array[7564] = 32'hFFFFFFF1;
    // rom_array[7565] = 32'h000053f9;
    // rom_array[7566] = 32'h00005401;
    // rom_array[7567] = 32'h00005409;
    // rom_array[7568] = 32'h00005411;
    // rom_array[7569] = 32'h00005419;
    // rom_array[7570] = 32'h00005421;
    // rom_array[7571] = 32'hFFFFFFF0;
    // rom_array[7572] = 32'hFFFFFFF0;
    // rom_array[7573] = 32'h00005429;
    // rom_array[7574] = 32'h00005431;
    // rom_array[7575] = 32'hFFFFFFF0;
    // rom_array[7576] = 32'hFFFFFFF0;
    // rom_array[7577] = 32'hFFFFFFF1;
    // rom_array[7578] = 32'hFFFFFFF1;
    // rom_array[7579] = 32'hFFFFFFF1;
    // rom_array[7580] = 32'hFFFFFFF1;
    // rom_array[7581] = 32'h00005439;
    // rom_array[7582] = 32'h00005441;
    // rom_array[7583] = 32'h00005449;
    // rom_array[7584] = 32'h00005451;
    // rom_array[7585] = 32'h00005459;
    // rom_array[7586] = 32'h00005461;
    // rom_array[7587] = 32'hFFFFFFF0;
    // rom_array[7588] = 32'hFFFFFFF0;
    // rom_array[7589] = 32'h00005469;
    // rom_array[7590] = 32'h00005471;
    // rom_array[7591] = 32'hFFFFFFF0;
    // rom_array[7592] = 32'hFFFFFFF0;
    // rom_array[7593] = 32'h00005479;
    // rom_array[7594] = 32'h00005481;
    // rom_array[7595] = 32'h00005489;
    // rom_array[7596] = 32'h00005491;
    // rom_array[7597] = 32'h00005499;
    // rom_array[7598] = 32'h000054a1;
    // rom_array[7599] = 32'h000054a9;
    // rom_array[7600] = 32'h000054b1;
    // rom_array[7601] = 32'h000054b9;
    // rom_array[7602] = 32'h000054c1;
    // rom_array[7603] = 32'h000054c9;
    // rom_array[7604] = 32'h000054d1;
    // rom_array[7605] = 32'h000054d9;
    // rom_array[7606] = 32'h000054e1;
    // rom_array[7607] = 32'h000054e9;
    // rom_array[7608] = 32'h000054f1;
    // rom_array[7609] = 32'h000054f9;
    // rom_array[7610] = 32'h00005501;
    // rom_array[7611] = 32'h00005509;
    // rom_array[7612] = 32'h00005511;
    // rom_array[7613] = 32'h00005519;
    // rom_array[7614] = 32'h00005521;
    // rom_array[7615] = 32'h00005529;
    // rom_array[7616] = 32'h00005531;
    // rom_array[7617] = 32'h00005539;
    // rom_array[7618] = 32'h00005541;
    // rom_array[7619] = 32'h00005549;
    // rom_array[7620] = 32'h00005551;
    // rom_array[7621] = 32'h00005559;
    // rom_array[7622] = 32'h00005561;
    // rom_array[7623] = 32'h00005569;
    // rom_array[7624] = 32'h00005571;
    // rom_array[7625] = 32'h00005579;
    // rom_array[7626] = 32'h00005581;
    // rom_array[7627] = 32'h00005589;
    // rom_array[7628] = 32'h00005591;
    // rom_array[7629] = 32'h00005599;
    // rom_array[7630] = 32'h000055a1;
    // rom_array[7631] = 32'h000055a9;
    // rom_array[7632] = 32'h000055b1;
    // rom_array[7633] = 32'h000055b9;
    // rom_array[7634] = 32'h000055c1;
    // rom_array[7635] = 32'hFFFFFFF0;
    // rom_array[7636] = 32'hFFFFFFF0;
    // rom_array[7637] = 32'h000055c9;
    // rom_array[7638] = 32'h000055d1;
    // rom_array[7639] = 32'h000055d9;
    // rom_array[7640] = 32'h000055e1;
    // rom_array[7641] = 32'h000055e9;
    // rom_array[7642] = 32'h000055f1;
    // rom_array[7643] = 32'h000055f9;
    // rom_array[7644] = 32'h00005601;
    // rom_array[7645] = 32'hFFFFFFF0;
    // rom_array[7646] = 32'hFFFFFFF0;
    // rom_array[7647] = 32'hFFFFFFF0;
    // rom_array[7648] = 32'hFFFFFFF0;
    // rom_array[7649] = 32'h00005609;
    // rom_array[7650] = 32'h00005611;
    // rom_array[7651] = 32'h00005619;
    // rom_array[7652] = 32'h00005621;
    // rom_array[7653] = 32'hFFFFFFF0;
    // rom_array[7654] = 32'hFFFFFFF0;
    // rom_array[7655] = 32'hFFFFFFF0;
    // rom_array[7656] = 32'hFFFFFFF0;
    // rom_array[7657] = 32'h00005629;
    // rom_array[7658] = 32'h00005631;
    // rom_array[7659] = 32'h00005639;
    // rom_array[7660] = 32'h00005641;
    // rom_array[7661] = 32'hFFFFFFF0;
    // rom_array[7662] = 32'hFFFFFFF0;
    // rom_array[7663] = 32'hFFFFFFF0;
    // rom_array[7664] = 32'hFFFFFFF0;
    // rom_array[7665] = 32'h00005649;
    // rom_array[7666] = 32'h00005651;
    // rom_array[7667] = 32'h00005659;
    // rom_array[7668] = 32'h00005661;
    // rom_array[7669] = 32'hFFFFFFF0;
    // rom_array[7670] = 32'hFFFFFFF0;
    // rom_array[7671] = 32'hFFFFFFF0;
    // rom_array[7672] = 32'hFFFFFFF0;
    // rom_array[7673] = 32'h00005669;
    // rom_array[7674] = 32'h00005671;
    // rom_array[7675] = 32'h00005679;
    // rom_array[7676] = 32'h00005681;
    // rom_array[7677] = 32'h00005689;
    // rom_array[7678] = 32'h00005691;
    // rom_array[7679] = 32'h00005699;
    // rom_array[7680] = 32'h000056a1;
    // rom_array[7681] = 32'h000056a9;
    // rom_array[7682] = 32'h000056b1;
    // rom_array[7683] = 32'h000056b9;
    // rom_array[7684] = 32'h000056c1;
    // rom_array[7685] = 32'hFFFFFFF0;
    // rom_array[7686] = 32'hFFFFFFF0;
    // rom_array[7687] = 32'hFFFFFFF0;
    // rom_array[7688] = 32'hFFFFFFF0;
    // rom_array[7689] = 32'h000056c9;
    // rom_array[7690] = 32'h000056d1;
    // rom_array[7691] = 32'h000056d9;
    // rom_array[7692] = 32'h000056e1;
    // rom_array[7693] = 32'hFFFFFFF1;
    // rom_array[7694] = 32'hFFFFFFF1;
    // rom_array[7695] = 32'h000056e9;
    // rom_array[7696] = 32'h000056f1;
    // rom_array[7697] = 32'hFFFFFFF1;
    // rom_array[7698] = 32'hFFFFFFF1;
    // rom_array[7699] = 32'h000056f9;
    // rom_array[7700] = 32'h00005701;
    // rom_array[7701] = 32'hFFFFFFF1;
    // rom_array[7702] = 32'hFFFFFFF1;
    // rom_array[7703] = 32'h00005709;
    // rom_array[7704] = 32'h00005711;
    // rom_array[7705] = 32'hFFFFFFF1;
    // rom_array[7706] = 32'hFFFFFFF1;
    // rom_array[7707] = 32'h00005719;
    // rom_array[7708] = 32'h00005721;
    // rom_array[7709] = 32'hFFFFFFF1;
    // rom_array[7710] = 32'hFFFFFFF1;
    // rom_array[7711] = 32'h00005729;
    // rom_array[7712] = 32'h00005731;
    // rom_array[7713] = 32'h00005739;
    // rom_array[7714] = 32'h00005741;
    // rom_array[7715] = 32'h00005749;
    // rom_array[7716] = 32'h00005751;
    // rom_array[7717] = 32'hFFFFFFF1;
    // rom_array[7718] = 32'hFFFFFFF1;
    // rom_array[7719] = 32'hFFFFFFF1;
    // rom_array[7720] = 32'hFFFFFFF1;
    // rom_array[7721] = 32'h00005759;
    // rom_array[7722] = 32'h00005761;
    // rom_array[7723] = 32'h00005769;
    // rom_array[7724] = 32'h00005771;
    // rom_array[7725] = 32'hFFFFFFF1;
    // rom_array[7726] = 32'hFFFFFFF1;
    // rom_array[7727] = 32'hFFFFFFF1;
    // rom_array[7728] = 32'hFFFFFFF1;
    // rom_array[7729] = 32'h00005779;
    // rom_array[7730] = 32'h00005781;
    // rom_array[7731] = 32'h00005789;
    // rom_array[7732] = 32'h00005791;
    // rom_array[7733] = 32'hFFFFFFF0;
    // rom_array[7734] = 32'hFFFFFFF0;
    // rom_array[7735] = 32'hFFFFFFF0;
    // rom_array[7736] = 32'hFFFFFFF0;
    // rom_array[7737] = 32'h00005799;
    // rom_array[7738] = 32'h000057a1;
    // rom_array[7739] = 32'h000057a9;
    // rom_array[7740] = 32'h000057b1;
    // rom_array[7741] = 32'hFFFFFFF0;
    // rom_array[7742] = 32'hFFFFFFF0;
    // rom_array[7743] = 32'hFFFFFFF0;
    // rom_array[7744] = 32'hFFFFFFF0;
    // rom_array[7745] = 32'h000057b9;
    // rom_array[7746] = 32'h000057c1;
    // rom_array[7747] = 32'h000057c9;
    // rom_array[7748] = 32'h000057d1;
    // rom_array[7749] = 32'hFFFFFFF1;
    // rom_array[7750] = 32'hFFFFFFF1;
    // rom_array[7751] = 32'hFFFFFFF1;
    // rom_array[7752] = 32'hFFFFFFF1;
    // rom_array[7753] = 32'h000057d9;
    // rom_array[7754] = 32'h000057e1;
    // rom_array[7755] = 32'h000057e9;
    // rom_array[7756] = 32'h000057f1;
    // rom_array[7757] = 32'hFFFFFFF1;
    // rom_array[7758] = 32'hFFFFFFF1;
    // rom_array[7759] = 32'hFFFFFFF1;
    // rom_array[7760] = 32'hFFFFFFF1;
    // rom_array[7761] = 32'h000057f9;
    // rom_array[7762] = 32'h00005801;
    // rom_array[7763] = 32'h00005809;
    // rom_array[7764] = 32'h00005811;
    // rom_array[7765] = 32'hFFFFFFF0;
    // rom_array[7766] = 32'hFFFFFFF0;
    // rom_array[7767] = 32'hFFFFFFF0;
    // rom_array[7768] = 32'hFFFFFFF0;
    // rom_array[7769] = 32'h00005819;
    // rom_array[7770] = 32'h00005821;
    // rom_array[7771] = 32'h00005829;
    // rom_array[7772] = 32'h00005831;
    // rom_array[7773] = 32'hFFFFFFF0;
    // rom_array[7774] = 32'hFFFFFFF0;
    // rom_array[7775] = 32'hFFFFFFF0;
    // rom_array[7776] = 32'hFFFFFFF0;
    // rom_array[7777] = 32'h00005839;
    // rom_array[7778] = 32'h00005841;
    // rom_array[7779] = 32'h00005849;
    // rom_array[7780] = 32'h00005851;
    // rom_array[7781] = 32'hFFFFFFF1;
    // rom_array[7782] = 32'hFFFFFFF1;
    // rom_array[7783] = 32'hFFFFFFF1;
    // rom_array[7784] = 32'hFFFFFFF1;
    // rom_array[7785] = 32'h00005859;
    // rom_array[7786] = 32'h00005861;
    // rom_array[7787] = 32'h00005869;
    // rom_array[7788] = 32'h00005871;
    // rom_array[7789] = 32'hFFFFFFF1;
    // rom_array[7790] = 32'hFFFFFFF1;
    // rom_array[7791] = 32'h00005879;
    // rom_array[7792] = 32'h00005881;
    // rom_array[7793] = 32'h00005889;
    // rom_array[7794] = 32'h00005891;
    // rom_array[7795] = 32'h00005899;
    // rom_array[7796] = 32'h000058a1;
    // rom_array[7797] = 32'hFFFFFFF0;
    // rom_array[7798] = 32'hFFFFFFF0;
    // rom_array[7799] = 32'hFFFFFFF0;
    // rom_array[7800] = 32'hFFFFFFF0;
    // rom_array[7801] = 32'h000058a9;
    // rom_array[7802] = 32'h000058b1;
    // rom_array[7803] = 32'h000058b9;
    // rom_array[7804] = 32'h000058c1;
    // rom_array[7805] = 32'hFFFFFFF1;
    // rom_array[7806] = 32'hFFFFFFF1;
    // rom_array[7807] = 32'h000058c9;
    // rom_array[7808] = 32'h000058d1;
    // rom_array[7809] = 32'hFFFFFFF1;
    // rom_array[7810] = 32'hFFFFFFF1;
    // rom_array[7811] = 32'h000058d9;
    // rom_array[7812] = 32'h000058e1;
    // rom_array[7813] = 32'hFFFFFFF1;
    // rom_array[7814] = 32'hFFFFFFF1;
    // rom_array[7815] = 32'h000058e9;
    // rom_array[7816] = 32'h000058f1;
    // rom_array[7817] = 32'hFFFFFFF1;
    // rom_array[7818] = 32'hFFFFFFF1;
    // rom_array[7819] = 32'h000058f9;
    // rom_array[7820] = 32'h00005901;
    // rom_array[7821] = 32'hFFFFFFF1;
    // rom_array[7822] = 32'hFFFFFFF1;
    // rom_array[7823] = 32'h00005909;
    // rom_array[7824] = 32'h00005911;
    // rom_array[7825] = 32'h00005919;
    // rom_array[7826] = 32'h00005921;
    // rom_array[7827] = 32'h00005929;
    // rom_array[7828] = 32'h00005931;
    // rom_array[7829] = 32'hFFFFFFF1;
    // rom_array[7830] = 32'hFFFFFFF1;
    // rom_array[7831] = 32'hFFFFFFF1;
    // rom_array[7832] = 32'hFFFFFFF1;
    // rom_array[7833] = 32'h00005939;
    // rom_array[7834] = 32'h00005941;
    // rom_array[7835] = 32'h00005949;
    // rom_array[7836] = 32'h00005951;
    // rom_array[7837] = 32'hFFFFFFF1;
    // rom_array[7838] = 32'hFFFFFFF1;
    // rom_array[7839] = 32'hFFFFFFF1;
    // rom_array[7840] = 32'hFFFFFFF1;
    // rom_array[7841] = 32'hFFFFFFF1;
    // rom_array[7842] = 32'hFFFFFFF1;
    // rom_array[7843] = 32'hFFFFFFF1;
    // rom_array[7844] = 32'hFFFFFFF1;
    // rom_array[7845] = 32'h00005959;
    // rom_array[7846] = 32'h00005961;
    // rom_array[7847] = 32'h00005969;
    // rom_array[7848] = 32'h00005971;
    // rom_array[7849] = 32'hFFFFFFF1;
    // rom_array[7850] = 32'hFFFFFFF1;
    // rom_array[7851] = 32'hFFFFFFF1;
    // rom_array[7852] = 32'hFFFFFFF1;
    // rom_array[7853] = 32'h00005979;
    // rom_array[7854] = 32'h00005981;
    // rom_array[7855] = 32'h00005989;
    // rom_array[7856] = 32'h00005991;
    // rom_array[7857] = 32'h00005999;
    // rom_array[7858] = 32'h000059a1;
    // rom_array[7859] = 32'h000059a9;
    // rom_array[7860] = 32'h000059b1;
    // rom_array[7861] = 32'hFFFFFFF1;
    // rom_array[7862] = 32'hFFFFFFF1;
    // rom_array[7863] = 32'hFFFFFFF1;
    // rom_array[7864] = 32'hFFFFFFF1;
    // rom_array[7865] = 32'h000059b9;
    // rom_array[7866] = 32'h000059c1;
    // rom_array[7867] = 32'h000059c9;
    // rom_array[7868] = 32'h000059d1;
    // rom_array[7869] = 32'hFFFFFFF1;
    // rom_array[7870] = 32'hFFFFFFF1;
    // rom_array[7871] = 32'hFFFFFFF1;
    // rom_array[7872] = 32'hFFFFFFF1;
    // rom_array[7873] = 32'hFFFFFFF1;
    // rom_array[7874] = 32'hFFFFFFF1;
    // rom_array[7875] = 32'hFFFFFFF1;
    // rom_array[7876] = 32'hFFFFFFF1;
    // rom_array[7877] = 32'h000059d9;
    // rom_array[7878] = 32'h000059e1;
    // rom_array[7879] = 32'h000059e9;
    // rom_array[7880] = 32'h000059f1;
    // rom_array[7881] = 32'hFFFFFFF1;
    // rom_array[7882] = 32'hFFFFFFF1;
    // rom_array[7883] = 32'hFFFFFFF1;
    // rom_array[7884] = 32'hFFFFFFF1;
    // rom_array[7885] = 32'h000059f9;
    // rom_array[7886] = 32'h00005a01;
    // rom_array[7887] = 32'h00005a09;
    // rom_array[7888] = 32'h00005a11;
    // rom_array[7889] = 32'h00005a19;
    // rom_array[7890] = 32'h00005a21;
    // rom_array[7891] = 32'h00005a29;
    // rom_array[7892] = 32'h00005a31;
    // rom_array[7893] = 32'hFFFFFFF0;
    // rom_array[7894] = 32'hFFFFFFF0;
    // rom_array[7895] = 32'hFFFFFFF0;
    // rom_array[7896] = 32'hFFFFFFF0;
    // rom_array[7897] = 32'h00005a39;
    // rom_array[7898] = 32'h00005a41;
    // rom_array[7899] = 32'h00005a49;
    // rom_array[7900] = 32'h00005a51;
    // rom_array[7901] = 32'hFFFFFFF0;
    // rom_array[7902] = 32'hFFFFFFF0;
    // rom_array[7903] = 32'hFFFFFFF0;
    // rom_array[7904] = 32'hFFFFFFF0;
    // rom_array[7905] = 32'h00005a59;
    // rom_array[7906] = 32'h00005a61;
    // rom_array[7907] = 32'h00005a69;
    // rom_array[7908] = 32'h00005a71;
    // rom_array[7909] = 32'hFFFFFFF0;
    // rom_array[7910] = 32'hFFFFFFF0;
    // rom_array[7911] = 32'hFFFFFFF0;
    // rom_array[7912] = 32'hFFFFFFF0;
    // rom_array[7913] = 32'h00005a79;
    // rom_array[7914] = 32'h00005a81;
    // rom_array[7915] = 32'h00005a89;
    // rom_array[7916] = 32'h00005a91;
    // rom_array[7917] = 32'hFFFFFFF0;
    // rom_array[7918] = 32'hFFFFFFF0;
    // rom_array[7919] = 32'hFFFFFFF0;
    // rom_array[7920] = 32'hFFFFFFF0;
    // rom_array[7921] = 32'h00005a99;
    // rom_array[7922] = 32'h00005aa1;
    // rom_array[7923] = 32'h00005aa9;
    // rom_array[7924] = 32'h00005ab1;
    // rom_array[7925] = 32'hFFFFFFF1;
    // rom_array[7926] = 32'hFFFFFFF1;
    // rom_array[7927] = 32'hFFFFFFF1;
    // rom_array[7928] = 32'hFFFFFFF1;
    // rom_array[7929] = 32'h00005ab9;
    // rom_array[7930] = 32'h00005ac1;
    // rom_array[7931] = 32'h00005ac9;
    // rom_array[7932] = 32'h00005ad1;
    // rom_array[7933] = 32'h00005ad9;
    // rom_array[7934] = 32'h00005ae1;
    // rom_array[7935] = 32'h00005ae9;
    // rom_array[7936] = 32'h00005af1;
    // rom_array[7937] = 32'hFFFFFFF1;
    // rom_array[7938] = 32'hFFFFFFF1;
    // rom_array[7939] = 32'hFFFFFFF1;
    // rom_array[7940] = 32'hFFFFFFF1;
    // rom_array[7941] = 32'h00005af9;
    // rom_array[7942] = 32'h00005b01;
    // rom_array[7943] = 32'h00005b09;
    // rom_array[7944] = 32'h00005b11;
    // rom_array[7945] = 32'h00005b19;
    // rom_array[7946] = 32'h00005b21;
    // rom_array[7947] = 32'h00005b29;
    // rom_array[7948] = 32'h00005b31;
    // rom_array[7949] = 32'h00005b39;
    // rom_array[7950] = 32'h00005b41;
    // rom_array[7951] = 32'h00005b49;
    // rom_array[7952] = 32'h00005b51;
    // rom_array[7953] = 32'h00005b59;
    // rom_array[7954] = 32'h00005b61;
    // rom_array[7955] = 32'h00005b69;
    // rom_array[7956] = 32'h00005b71;
    // rom_array[7957] = 32'hFFFFFFF0;
    // rom_array[7958] = 32'hFFFFFFF0;
    // rom_array[7959] = 32'hFFFFFFF0;
    // rom_array[7960] = 32'hFFFFFFF0;
    // rom_array[7961] = 32'h00005b79;
    // rom_array[7962] = 32'h00005b81;
    // rom_array[7963] = 32'hFFFFFFF0;
    // rom_array[7964] = 32'hFFFFFFF0;
    // rom_array[7965] = 32'hFFFFFFF0;
    // rom_array[7966] = 32'hFFFFFFF0;
    // rom_array[7967] = 32'hFFFFFFF0;
    // rom_array[7968] = 32'hFFFFFFF0;
    // rom_array[7969] = 32'h00005b89;
    // rom_array[7970] = 32'h00005b91;
    // rom_array[7971] = 32'h00005b99;
    // rom_array[7972] = 32'h00005ba1;
    // rom_array[7973] = 32'hFFFFFFF1;
    // rom_array[7974] = 32'hFFFFFFF1;
    // rom_array[7975] = 32'hFFFFFFF1;
    // rom_array[7976] = 32'hFFFFFFF1;
    // rom_array[7977] = 32'h00005ba9;
    // rom_array[7978] = 32'h00005bb1;
    // rom_array[7979] = 32'h00005bb9;
    // rom_array[7980] = 32'h00005bc1;
    // rom_array[7981] = 32'hFFFFFFF1;
    // rom_array[7982] = 32'hFFFFFFF1;
    // rom_array[7983] = 32'hFFFFFFF1;
    // rom_array[7984] = 32'hFFFFFFF1;
    // rom_array[7985] = 32'h00005bc9;
    // rom_array[7986] = 32'h00005bd1;
    // rom_array[7987] = 32'h00005bd9;
    // rom_array[7988] = 32'h00005be1;
    // rom_array[7989] = 32'hFFFFFFF1;
    // rom_array[7990] = 32'hFFFFFFF1;
    // rom_array[7991] = 32'hFFFFFFF1;
    // rom_array[7992] = 32'hFFFFFFF1;
    // rom_array[7993] = 32'h00005be9;
    // rom_array[7994] = 32'h00005bf1;
    // rom_array[7995] = 32'h00005bf9;
    // rom_array[7996] = 32'h00005c01;
    // rom_array[7997] = 32'hFFFFFFF1;
    // rom_array[7998] = 32'hFFFFFFF1;
    // rom_array[7999] = 32'hFFFFFFF1;
    // rom_array[8000] = 32'hFFFFFFF1;
    // rom_array[8001] = 32'h00005c09;
    // rom_array[8002] = 32'h00005c11;
    // rom_array[8003] = 32'h00005c19;
    // rom_array[8004] = 32'h00005c21;
    // rom_array[8005] = 32'h00005c29;
    // rom_array[8006] = 32'h00005c31;
    // rom_array[8007] = 32'hFFFFFFF0;
    // rom_array[8008] = 32'hFFFFFFF0;
    // rom_array[8009] = 32'h00005c39;
    // rom_array[8010] = 32'h00005c41;
    // rom_array[8011] = 32'h00005c49;
    // rom_array[8012] = 32'h00005c51;
    // rom_array[8013] = 32'hFFFFFFF0;
    // rom_array[8014] = 32'hFFFFFFF0;
    // rom_array[8015] = 32'hFFFFFFF0;
    // rom_array[8016] = 32'hFFFFFFF0;
    // rom_array[8017] = 32'h00005c59;
    // rom_array[8018] = 32'h00005c61;
    // rom_array[8019] = 32'hFFFFFFF0;
    // rom_array[8020] = 32'hFFFFFFF0;
    // rom_array[8021] = 32'h00005c69;
    // rom_array[8022] = 32'h00005c71;
    // rom_array[8023] = 32'hFFFFFFF0;
    // rom_array[8024] = 32'hFFFFFFF0;
    // rom_array[8025] = 32'h00005c79;
    // rom_array[8026] = 32'h00005c81;
    // rom_array[8027] = 32'h00005c89;
    // rom_array[8028] = 32'h00005c91;
    // rom_array[8029] = 32'hFFFFFFF0;
    // rom_array[8030] = 32'hFFFFFFF0;
    // rom_array[8031] = 32'hFFFFFFF0;
    // rom_array[8032] = 32'hFFFFFFF0;
    // rom_array[8033] = 32'h00005c99;
    // rom_array[8034] = 32'h00005ca1;
    // rom_array[8035] = 32'h00005ca9;
    // rom_array[8036] = 32'h00005cb1;
    // rom_array[8037] = 32'h00005cb9;
    // rom_array[8038] = 32'h00005cc1;
    // rom_array[8039] = 32'hFFFFFFF1;
    // rom_array[8040] = 32'hFFFFFFF1;
    // rom_array[8041] = 32'h00005cc9;
    // rom_array[8042] = 32'h00005cd1;
    // rom_array[8043] = 32'hFFFFFFF1;
    // rom_array[8044] = 32'hFFFFFFF1;
    // rom_array[8045] = 32'h00005cd9;
    // rom_array[8046] = 32'h00005ce1;
    // rom_array[8047] = 32'hFFFFFFF1;
    // rom_array[8048] = 32'hFFFFFFF1;
    // rom_array[8049] = 32'h00005ce9;
    // rom_array[8050] = 32'h00005cf1;
    // rom_array[8051] = 32'h00005cf9;
    // rom_array[8052] = 32'h00005d01;
    // rom_array[8053] = 32'hFFFFFFF1;
    // rom_array[8054] = 32'hFFFFFFF1;
    // rom_array[8055] = 32'hFFFFFFF1;
    // rom_array[8056] = 32'hFFFFFFF1;
    // rom_array[8057] = 32'h00005d09;
    // rom_array[8058] = 32'h00005d11;
    // rom_array[8059] = 32'hFFFFFFF0;
    // rom_array[8060] = 32'hFFFFFFF0;
    // rom_array[8061] = 32'h00005d19;
    // rom_array[8062] = 32'h00005d21;
    // rom_array[8063] = 32'hFFFFFFF0;
    // rom_array[8064] = 32'hFFFFFFF0;
    // rom_array[8065] = 32'h00005d29;
    // rom_array[8066] = 32'h00005d31;
    // rom_array[8067] = 32'hFFFFFFF0;
    // rom_array[8068] = 32'hFFFFFFF0;
    // rom_array[8069] = 32'h00005d39;
    // rom_array[8070] = 32'h00005d41;
    // rom_array[8071] = 32'hFFFFFFF0;
    // rom_array[8072] = 32'hFFFFFFF0;
    // rom_array[8073] = 32'h00005d49;
    // rom_array[8074] = 32'h00005d51;
    // rom_array[8075] = 32'h00005d59;
    // rom_array[8076] = 32'h00005d61;
    // rom_array[8077] = 32'hFFFFFFF1;
    // rom_array[8078] = 32'hFFFFFFF1;
    // rom_array[8079] = 32'hFFFFFFF1;
    // rom_array[8080] = 32'hFFFFFFF1;
    // rom_array[8081] = 32'h00005d69;
    // rom_array[8082] = 32'h00005d71;
    // rom_array[8083] = 32'hFFFFFFF0;
    // rom_array[8084] = 32'hFFFFFFF0;
    // rom_array[8085] = 32'h00005d79;
    // rom_array[8086] = 32'h00005d81;
    // rom_array[8087] = 32'hFFFFFFF0;
    // rom_array[8088] = 32'hFFFFFFF0;
    // rom_array[8089] = 32'h00005d89;
    // rom_array[8090] = 32'h00005d91;
    // rom_array[8091] = 32'hFFFFFFF0;
    // rom_array[8092] = 32'hFFFFFFF0;
    // rom_array[8093] = 32'h00005d99;
    // rom_array[8094] = 32'h00005da1;
    // rom_array[8095] = 32'hFFFFFFF0;
    // rom_array[8096] = 32'hFFFFFFF0;
    // rom_array[8097] = 32'h00005da9;
    // rom_array[8098] = 32'h00005db1;
    // rom_array[8099] = 32'hFFFFFFF0;
    // rom_array[8100] = 32'hFFFFFFF0;
    // rom_array[8101] = 32'h00005db9;
    // rom_array[8102] = 32'h00005dc1;
    // rom_array[8103] = 32'hFFFFFFF0;
    // rom_array[8104] = 32'hFFFFFFF0;
    // rom_array[8105] = 32'h00005dc9;
    // rom_array[8106] = 32'h00005dd1;
    // rom_array[8107] = 32'hFFFFFFF0;
    // rom_array[8108] = 32'hFFFFFFF0;
    // rom_array[8109] = 32'h00005dd9;
    // rom_array[8110] = 32'h00005de1;
    // rom_array[8111] = 32'h00005de9;
    // rom_array[8112] = 32'h00005df1;
    // rom_array[8113] = 32'hFFFFFFF0;
    // rom_array[8114] = 32'hFFFFFFF0;
    // rom_array[8115] = 32'hFFFFFFF0;
    // rom_array[8116] = 32'hFFFFFFF0;
    // rom_array[8117] = 32'h00005df9;
    // rom_array[8118] = 32'h00005e01;
    // rom_array[8119] = 32'h00005e09;
    // rom_array[8120] = 32'h00005e11;
    // rom_array[8121] = 32'h00005e19;
    // rom_array[8122] = 32'h00005e21;
    // rom_array[8123] = 32'hFFFFFFF1;
    // rom_array[8124] = 32'hFFFFFFF1;
    // rom_array[8125] = 32'h00005e29;
    // rom_array[8126] = 32'h00005e31;
    // rom_array[8127] = 32'hFFFFFFF1;
    // rom_array[8128] = 32'hFFFFFFF1;
    // rom_array[8129] = 32'hFFFFFFF0;
    // rom_array[8130] = 32'hFFFFFFF0;
    // rom_array[8131] = 32'hFFFFFFF0;
    // rom_array[8132] = 32'hFFFFFFF0;
    // rom_array[8133] = 32'h00005e39;
    // rom_array[8134] = 32'h00005e41;
    // rom_array[8135] = 32'h00005e49;
    // rom_array[8136] = 32'h00005e51;
    // rom_array[8137] = 32'h00005e59;
    // rom_array[8138] = 32'h00005e61;
    // rom_array[8139] = 32'hFFFFFFF1;
    // rom_array[8140] = 32'hFFFFFFF1;
    // rom_array[8141] = 32'h00005e69;
    // rom_array[8142] = 32'h00005e71;
    // rom_array[8143] = 32'h00005e79;
    // rom_array[8144] = 32'h00005e81;
    // rom_array[8145] = 32'h00005e89;
    // rom_array[8146] = 32'h00005e91;
    // rom_array[8147] = 32'hFFFFFFF0;
    // rom_array[8148] = 32'hFFFFFFF0;
    // rom_array[8149] = 32'hFFFFFFF0;
    // rom_array[8150] = 32'hFFFFFFF0;
    // rom_array[8151] = 32'hFFFFFFF0;
    // rom_array[8152] = 32'hFFFFFFF0;
    // rom_array[8153] = 32'hFFFFFFF1;
    // rom_array[8154] = 32'hFFFFFFF1;
    // rom_array[8155] = 32'hFFFFFFF1;
    // rom_array[8156] = 32'hFFFFFFF1;
    // rom_array[8157] = 32'h00005e99;
    // rom_array[8158] = 32'h00005ea1;
    // rom_array[8159] = 32'h00005ea9;
    // rom_array[8160] = 32'h00005eb1;
    // rom_array[8161] = 32'hFFFFFFF1;
    // rom_array[8162] = 32'hFFFFFFF1;
    // rom_array[8163] = 32'hFFFFFFF1;
    // rom_array[8164] = 32'hFFFFFFF1;
    // rom_array[8165] = 32'h00005eb9;
    // rom_array[8166] = 32'h00005ec1;
    // rom_array[8167] = 32'h00005ec9;
    // rom_array[8168] = 32'h00005ed1;
    // rom_array[8169] = 32'h00005ed9;
    // rom_array[8170] = 32'h00005ee1;
    // rom_array[8171] = 32'h00005ee9;
    // rom_array[8172] = 32'h00005ef1;
    // rom_array[8173] = 32'hFFFFFFF1;
    // rom_array[8174] = 32'hFFFFFFF1;
    // rom_array[8175] = 32'h00005ef9;
    // rom_array[8176] = 32'h00005f01;
    // rom_array[8177] = 32'hFFFFFFF1;
    // rom_array[8178] = 32'hFFFFFFF1;
    // rom_array[8179] = 32'hFFFFFFF1;
    // rom_array[8180] = 32'hFFFFFFF1;
    // rom_array[8181] = 32'h00005f09;
    // rom_array[8182] = 32'h00005f11;
    // rom_array[8183] = 32'h00005f19;
    // rom_array[8184] = 32'h00005f21;
    // rom_array[8185] = 32'hFFFFFFF1;
    // rom_array[8186] = 32'hFFFFFFF1;
    // rom_array[8187] = 32'h00005f29;
    // rom_array[8188] = 32'h00005f31;
    // rom_array[8189] = 32'h00005f39;
    // rom_array[8190] = 32'h00005f41;
    // rom_array[8191] = 32'h00005f49;
    // rom_array[8192] = 32'h00005f51;
    // rom_array[8193] = 32'h00005f59;
    // rom_array[8194] = 32'h00005f61;
    // rom_array[8195] = 32'hFFFFFFF0;
    // rom_array[8196] = 32'hFFFFFFF0;
    // rom_array[8197] = 32'h00005f69;
    // rom_array[8198] = 32'h00005f71;
    // rom_array[8199] = 32'hFFFFFFF0;
    // rom_array[8200] = 32'hFFFFFFF0;
    // rom_array[8201] = 32'h00005f79;
    // rom_array[8202] = 32'h00005f81;
    // rom_array[8203] = 32'hFFFFFFF0;
    // rom_array[8204] = 32'hFFFFFFF0;
    // rom_array[8205] = 32'h00005f89;
    // rom_array[8206] = 32'h00005f91;
    // rom_array[8207] = 32'hFFFFFFF0;
    // rom_array[8208] = 32'hFFFFFFF0;
    // rom_array[8209] = 32'h00005f99;
    // rom_array[8210] = 32'h00005fa1;
    // rom_array[8211] = 32'h00005fa9;
    // rom_array[8212] = 32'h00005fb1;
    // rom_array[8213] = 32'hFFFFFFF0;
    // rom_array[8214] = 32'hFFFFFFF0;
    // rom_array[8215] = 32'hFFFFFFF0;
    // rom_array[8216] = 32'hFFFFFFF0;
    // rom_array[8217] = 32'h00005fb9;
    // rom_array[8218] = 32'h00005fc1;
    // rom_array[8219] = 32'hFFFFFFF0;
    // rom_array[8220] = 32'hFFFFFFF0;
    // rom_array[8221] = 32'hFFFFFFF0;
    // rom_array[8222] = 32'hFFFFFFF0;
    // rom_array[8223] = 32'hFFFFFFF0;
    // rom_array[8224] = 32'hFFFFFFF0;
    // rom_array[8225] = 32'h00005fc9;
    // rom_array[8226] = 32'h00005fd1;
    // rom_array[8227] = 32'h00005fd9;
    // rom_array[8228] = 32'h00005fe1;
    // rom_array[8229] = 32'hFFFFFFF1;
    // rom_array[8230] = 32'hFFFFFFF1;
    // rom_array[8231] = 32'hFFFFFFF1;
    // rom_array[8232] = 32'hFFFFFFF1;
    // rom_array[8233] = 32'h00005fe9;
    // rom_array[8234] = 32'h00005ff1;
    // rom_array[8235] = 32'h00005ff9;
    // rom_array[8236] = 32'h00006001;
    // rom_array[8237] = 32'hFFFFFFF1;
    // rom_array[8238] = 32'hFFFFFFF1;
    // rom_array[8239] = 32'hFFFFFFF1;
    // rom_array[8240] = 32'hFFFFFFF1;
    // rom_array[8241] = 32'h00006009;
    // rom_array[8242] = 32'h00006011;
    // rom_array[8243] = 32'h00006019;
    // rom_array[8244] = 32'h00006021;
    // rom_array[8245] = 32'hFFFFFFF1;
    // rom_array[8246] = 32'hFFFFFFF1;
    // rom_array[8247] = 32'hFFFFFFF1;
    // rom_array[8248] = 32'hFFFFFFF1;
    // rom_array[8249] = 32'h00006029;
    // rom_array[8250] = 32'h00006031;
    // rom_array[8251] = 32'h00006039;
    // rom_array[8252] = 32'h00006041;
    // rom_array[8253] = 32'hFFFFFFF1;
    // rom_array[8254] = 32'hFFFFFFF1;
    // rom_array[8255] = 32'hFFFFFFF1;
    // rom_array[8256] = 32'hFFFFFFF1;
    // rom_array[8257] = 32'h00006049;
    // rom_array[8258] = 32'h00006051;
    // rom_array[8259] = 32'h00006059;
    // rom_array[8260] = 32'h00006061;
    // rom_array[8261] = 32'hFFFFFFF1;
    // rom_array[8262] = 32'hFFFFFFF1;
    // rom_array[8263] = 32'h00006069;
    // rom_array[8264] = 32'h00006071;
    // rom_array[8265] = 32'h00006079;
    // rom_array[8266] = 32'h00006081;
    // rom_array[8267] = 32'h00006089;
    // rom_array[8268] = 32'h00006091;
    // rom_array[8269] = 32'hFFFFFFF0;
    // rom_array[8270] = 32'hFFFFFFF0;
    // rom_array[8271] = 32'hFFFFFFF0;
    // rom_array[8272] = 32'hFFFFFFF0;
    // rom_array[8273] = 32'h00006099;
    // rom_array[8274] = 32'h000060a1;
    // rom_array[8275] = 32'h000060a9;
    // rom_array[8276] = 32'h000060b1;
    // rom_array[8277] = 32'hFFFFFFF0;
    // rom_array[8278] = 32'hFFFFFFF0;
    // rom_array[8279] = 32'hFFFFFFF0;
    // rom_array[8280] = 32'hFFFFFFF0;
    // rom_array[8281] = 32'h000060b9;
    // rom_array[8282] = 32'h000060c1;
    // rom_array[8283] = 32'h000060c9;
    // rom_array[8284] = 32'h000060d1;
    // rom_array[8285] = 32'h000060d9;
    // rom_array[8286] = 32'h000060e1;
    // rom_array[8287] = 32'hFFFFFFF1;
    // rom_array[8288] = 32'hFFFFFFF1;
    // rom_array[8289] = 32'h000060e9;
    // rom_array[8290] = 32'h000060f1;
    // rom_array[8291] = 32'h000060f9;
    // rom_array[8292] = 32'h00006101;
    // rom_array[8293] = 32'hFFFFFFF1;
    // rom_array[8294] = 32'hFFFFFFF1;
    // rom_array[8295] = 32'hFFFFFFF1;
    // rom_array[8296] = 32'hFFFFFFF1;
    // rom_array[8297] = 32'h00006109;
    // rom_array[8298] = 32'h00006111;
    // rom_array[8299] = 32'hFFFFFFF0;
    // rom_array[8300] = 32'hFFFFFFF0;
    // rom_array[8301] = 32'h00006119;
    // rom_array[8302] = 32'h00006121;
    // rom_array[8303] = 32'hFFFFFFF0;
    // rom_array[8304] = 32'hFFFFFFF0;
    // rom_array[8305] = 32'h00006129;
    // rom_array[8306] = 32'h00006131;
    // rom_array[8307] = 32'hFFFFFFF0;
    // rom_array[8308] = 32'hFFFFFFF0;
    // rom_array[8309] = 32'h00006139;
    // rom_array[8310] = 32'h00006141;
    // rom_array[8311] = 32'hFFFFFFF0;
    // rom_array[8312] = 32'hFFFFFFF0;
    // rom_array[8313] = 32'h00006149;
    // rom_array[8314] = 32'h00006151;
    // rom_array[8315] = 32'h00006159;
    // rom_array[8316] = 32'h00006161;
    // rom_array[8317] = 32'hFFFFFFF1;
    // rom_array[8318] = 32'hFFFFFFF1;
    // rom_array[8319] = 32'hFFFFFFF1;
    // rom_array[8320] = 32'hFFFFFFF1;
    // rom_array[8321] = 32'h00006169;
    // rom_array[8322] = 32'h00006171;
    // rom_array[8323] = 32'hFFFFFFF0;
    // rom_array[8324] = 32'hFFFFFFF0;
    // rom_array[8325] = 32'h00006179;
    // rom_array[8326] = 32'h00006181;
    // rom_array[8327] = 32'hFFFFFFF0;
    // rom_array[8328] = 32'hFFFFFFF0;
    // rom_array[8329] = 32'hFFFFFFF1;
    // rom_array[8330] = 32'hFFFFFFF1;
    // rom_array[8331] = 32'h00006189;
    // rom_array[8332] = 32'h00006191;
    // rom_array[8333] = 32'hFFFFFFF1;
    // rom_array[8334] = 32'hFFFFFFF1;
    // rom_array[8335] = 32'h00006199;
    // rom_array[8336] = 32'h000061a1;
    // rom_array[8337] = 32'hFFFFFFF1;
    // rom_array[8338] = 32'hFFFFFFF1;
    // rom_array[8339] = 32'h000061a9;
    // rom_array[8340] = 32'h000061b1;
    // rom_array[8341] = 32'hFFFFFFF1;
    // rom_array[8342] = 32'hFFFFFFF1;
    // rom_array[8343] = 32'h000061b9;
    // rom_array[8344] = 32'h000061c1;
    // rom_array[8345] = 32'h000061c9;
    // rom_array[8346] = 32'h000061d1;
    // rom_array[8347] = 32'hFFFFFFF1;
    // rom_array[8348] = 32'hFFFFFFF1;
    // rom_array[8349] = 32'h000061d9;
    // rom_array[8350] = 32'h000061e1;
    // rom_array[8351] = 32'hFFFFFFF1;
    // rom_array[8352] = 32'hFFFFFFF1;
    // rom_array[8353] = 32'h000061e9;
    // rom_array[8354] = 32'h000061f1;
    // rom_array[8355] = 32'hFFFFFFF1;
    // rom_array[8356] = 32'hFFFFFFF1;
    // rom_array[8357] = 32'h000061f9;
    // rom_array[8358] = 32'h00006201;
    // rom_array[8359] = 32'hFFFFFFF1;
    // rom_array[8360] = 32'hFFFFFFF1;
    // rom_array[8361] = 32'hFFFFFFF1;
    // rom_array[8362] = 32'hFFFFFFF1;
    // rom_array[8363] = 32'h00006209;
    // rom_array[8364] = 32'h00006211;
    // rom_array[8365] = 32'hFFFFFFF1;
    // rom_array[8366] = 32'hFFFFFFF1;
    // rom_array[8367] = 32'h00006219;
    // rom_array[8368] = 32'h00006221;
    // rom_array[8369] = 32'hFFFFFFF1;
    // rom_array[8370] = 32'hFFFFFFF1;
    // rom_array[8371] = 32'h00006229;
    // rom_array[8372] = 32'h00006231;
    // rom_array[8373] = 32'hFFFFFFF1;
    // rom_array[8374] = 32'hFFFFFFF1;
    // rom_array[8375] = 32'h00006239;
    // rom_array[8376] = 32'h00006241;
    // rom_array[8377] = 32'h00006249;
    // rom_array[8378] = 32'h00006251;
    // rom_array[8379] = 32'hFFFFFFF1;
    // rom_array[8380] = 32'hFFFFFFF1;
    // rom_array[8381] = 32'h00006259;
    // rom_array[8382] = 32'h00006261;
    // rom_array[8383] = 32'hFFFFFFF1;
    // rom_array[8384] = 32'hFFFFFFF1;
    // rom_array[8385] = 32'h00006269;
    // rom_array[8386] = 32'h00006271;
    // rom_array[8387] = 32'hFFFFFFF1;
    // rom_array[8388] = 32'hFFFFFFF1;
    // rom_array[8389] = 32'h00006279;
    // rom_array[8390] = 32'h00006281;
    // rom_array[8391] = 32'hFFFFFFF1;
    // rom_array[8392] = 32'hFFFFFFF1;
    // rom_array[8393] = 32'h00006289;
    // rom_array[8394] = 32'h00006291;
    // rom_array[8395] = 32'hFFFFFFF0;
    // rom_array[8396] = 32'hFFFFFFF0;
    // rom_array[8397] = 32'h00006299;
    // rom_array[8398] = 32'h000062a1;
    // rom_array[8399] = 32'hFFFFFFF0;
    // rom_array[8400] = 32'hFFFFFFF0;
    // rom_array[8401] = 32'h000062a9;
    // rom_array[8402] = 32'h000062b1;
    // rom_array[8403] = 32'hFFFFFFF0;
    // rom_array[8404] = 32'hFFFFFFF0;
    // rom_array[8405] = 32'h000062b9;
    // rom_array[8406] = 32'h000062c1;
    // rom_array[8407] = 32'hFFFFFFF0;
    // rom_array[8408] = 32'hFFFFFFF0;
    // rom_array[8409] = 32'h000062c9;
    // rom_array[8410] = 32'h000062d1;
    // rom_array[8411] = 32'hFFFFFFF0;
    // rom_array[8412] = 32'hFFFFFFF0;
    // rom_array[8413] = 32'h000062d9;
    // rom_array[8414] = 32'h000062e1;
    // rom_array[8415] = 32'hFFFFFFF0;
    // rom_array[8416] = 32'hFFFFFFF0;
    // rom_array[8417] = 32'h000062e9;
    // rom_array[8418] = 32'h000062f1;
    // rom_array[8419] = 32'hFFFFFFF0;
    // rom_array[8420] = 32'hFFFFFFF0;
    // rom_array[8421] = 32'h000062f9;
    // rom_array[8422] = 32'h00006301;
    // rom_array[8423] = 32'hFFFFFFF0;
    // rom_array[8424] = 32'hFFFFFFF0;
    // rom_array[8425] = 32'hFFFFFFF0;
    // rom_array[8426] = 32'hFFFFFFF0;
    // rom_array[8427] = 32'hFFFFFFF0;
    // rom_array[8428] = 32'hFFFFFFF0;
    // rom_array[8429] = 32'h00006309;
    // rom_array[8430] = 32'h00006311;
    // rom_array[8431] = 32'h00006319;
    // rom_array[8432] = 32'h00006321;
    // rom_array[8433] = 32'h00006329;
    // rom_array[8434] = 32'h00006331;
    // rom_array[8435] = 32'hFFFFFFF1;
    // rom_array[8436] = 32'hFFFFFFF1;
    // rom_array[8437] = 32'h00006339;
    // rom_array[8438] = 32'h00006341;
    // rom_array[8439] = 32'hFFFFFFF1;
    // rom_array[8440] = 32'hFFFFFFF1;
    // rom_array[8441] = 32'hFFFFFFF0;
    // rom_array[8442] = 32'hFFFFFFF0;
    // rom_array[8443] = 32'hFFFFFFF0;
    // rom_array[8444] = 32'hFFFFFFF0;
    // rom_array[8445] = 32'h00006349;
    // rom_array[8446] = 32'h00006351;
    // rom_array[8447] = 32'h00006359;
    // rom_array[8448] = 32'h00006361;
    // rom_array[8449] = 32'hFFFFFFF0;
    // rom_array[8450] = 32'hFFFFFFF0;
    // rom_array[8451] = 32'hFFFFFFF0;
    // rom_array[8452] = 32'hFFFFFFF0;
    // rom_array[8453] = 32'h00006369;
    // rom_array[8454] = 32'h00006371;
    // rom_array[8455] = 32'hFFFFFFF0;
    // rom_array[8456] = 32'hFFFFFFF0;
    // rom_array[8457] = 32'h00006379;
    // rom_array[8458] = 32'h00006381;
    // rom_array[8459] = 32'hFFFFFFF0;
    // rom_array[8460] = 32'hFFFFFFF0;
    // rom_array[8461] = 32'h00006389;
    // rom_array[8462] = 32'h00006391;
    // rom_array[8463] = 32'hFFFFFFF0;
    // rom_array[8464] = 32'hFFFFFFF0;
    // rom_array[8465] = 32'h00006399;
    // rom_array[8466] = 32'h000063a1;
    // rom_array[8467] = 32'h000063a9;
    // rom_array[8468] = 32'h000063b1;
    // rom_array[8469] = 32'hFFFFFFF1;
    // rom_array[8470] = 32'hFFFFFFF1;
    // rom_array[8471] = 32'hFFFFFFF1;
    // rom_array[8472] = 32'hFFFFFFF1;
    // rom_array[8473] = 32'h000063b9;
    // rom_array[8474] = 32'h000063c1;
    // rom_array[8475] = 32'h000063c9;
    // rom_array[8476] = 32'h000063d1;
    // rom_array[8477] = 32'hFFFFFFF1;
    // rom_array[8478] = 32'hFFFFFFF1;
    // rom_array[8479] = 32'hFFFFFFF1;
    // rom_array[8480] = 32'hFFFFFFF1;
    // rom_array[8481] = 32'h000063d9;
    // rom_array[8482] = 32'h000063e1;
    // rom_array[8483] = 32'hFFFFFFF1;
    // rom_array[8484] = 32'hFFFFFFF1;
    // rom_array[8485] = 32'h000063e9;
    // rom_array[8486] = 32'h000063f1;
    // rom_array[8487] = 32'hFFFFFFF1;
    // rom_array[8488] = 32'hFFFFFFF1;
    // rom_array[8489] = 32'h000063f9;
    // rom_array[8490] = 32'h00006401;
    // rom_array[8491] = 32'h00006409;
    // rom_array[8492] = 32'h00006411;
    // rom_array[8493] = 32'hFFFFFFF1;
    // rom_array[8494] = 32'hFFFFFFF1;
    // rom_array[8495] = 32'hFFFFFFF1;
    // rom_array[8496] = 32'hFFFFFFF1;
    // rom_array[8497] = 32'h00006419;
    // rom_array[8498] = 32'h00006421;
    // rom_array[8499] = 32'hFFFFFFF1;
    // rom_array[8500] = 32'hFFFFFFF1;
    // rom_array[8501] = 32'h00006429;
    // rom_array[8502] = 32'h00006431;
    // rom_array[8503] = 32'hFFFFFFF1;
    // rom_array[8504] = 32'hFFFFFFF1;
    // rom_array[8505] = 32'h00006439;
    // rom_array[8506] = 32'h00006441;
    // rom_array[8507] = 32'h00006449;
    // rom_array[8508] = 32'h00006451;
    // rom_array[8509] = 32'hFFFFFFF0;
    // rom_array[8510] = 32'hFFFFFFF0;
    // rom_array[8511] = 32'hFFFFFFF0;
    // rom_array[8512] = 32'hFFFFFFF0;
    // rom_array[8513] = 32'h00006459;
    // rom_array[8514] = 32'h00006461;
    // rom_array[8515] = 32'h00006469;
    // rom_array[8516] = 32'h00006471;
    // rom_array[8517] = 32'hFFFFFFF0;
    // rom_array[8518] = 32'hFFFFFFF0;
    // rom_array[8519] = 32'hFFFFFFF0;
    // rom_array[8520] = 32'hFFFFFFF0;
    // rom_array[8521] = 32'h00006479;
    // rom_array[8522] = 32'h00006481;
    // rom_array[8523] = 32'hFFFFFFF1;
    // rom_array[8524] = 32'hFFFFFFF1;
    // rom_array[8525] = 32'h00006489;
    // rom_array[8526] = 32'h00006491;
    // rom_array[8527] = 32'hFFFFFFF1;
    // rom_array[8528] = 32'hFFFFFFF1;
    // rom_array[8529] = 32'h00006499;
    // rom_array[8530] = 32'h000064a1;
    // rom_array[8531] = 32'h000064a9;
    // rom_array[8532] = 32'h000064b1;
    // rom_array[8533] = 32'hFFFFFFF0;
    // rom_array[8534] = 32'hFFFFFFF0;
    // rom_array[8535] = 32'hFFFFFFF0;
    // rom_array[8536] = 32'hFFFFFFF0;
    // rom_array[8537] = 32'h000064b9;
    // rom_array[8538] = 32'h000064c1;
    // rom_array[8539] = 32'hFFFFFFF1;
    // rom_array[8540] = 32'hFFFFFFF1;
    // rom_array[8541] = 32'h000064c9;
    // rom_array[8542] = 32'h000064d1;
    // rom_array[8543] = 32'hFFFFFFF1;
    // rom_array[8544] = 32'hFFFFFFF1;
    // rom_array[8545] = 32'h000064d9;
    // rom_array[8546] = 32'h000064e1;
    // rom_array[8547] = 32'hFFFFFFF0;
    // rom_array[8548] = 32'hFFFFFFF0;
    // rom_array[8549] = 32'h000064e9;
    // rom_array[8550] = 32'h000064f1;
    // rom_array[8551] = 32'hFFFFFFF0;
    // rom_array[8552] = 32'hFFFFFFF0;
    // rom_array[8553] = 32'h000064f9;
    // rom_array[8554] = 32'h00006501;
    // rom_array[8555] = 32'hFFFFFFF0;
    // rom_array[8556] = 32'hFFFFFFF0;
    // rom_array[8557] = 32'h00006509;
    // rom_array[8558] = 32'h00006511;
    // rom_array[8559] = 32'hFFFFFFF0;
    // rom_array[8560] = 32'hFFFFFFF0;
    // rom_array[8561] = 32'h00006519;
    // rom_array[8562] = 32'h00006521;
    // rom_array[8563] = 32'hFFFFFFF0;
    // rom_array[8564] = 32'hFFFFFFF0;
    // rom_array[8565] = 32'h00006529;
    // rom_array[8566] = 32'h00006531;
    // rom_array[8567] = 32'hFFFFFFF0;
    // rom_array[8568] = 32'hFFFFFFF0;
    // rom_array[8569] = 32'h00006539;
    // rom_array[8570] = 32'h00006541;
    // rom_array[8571] = 32'hFFFFFFF0;
    // rom_array[8572] = 32'hFFFFFFF0;
    // rom_array[8573] = 32'h00006549;
    // rom_array[8574] = 32'h00006551;
    // rom_array[8575] = 32'hFFFFFFF0;
    // rom_array[8576] = 32'hFFFFFFF0;
    // rom_array[8577] = 32'h00006559;
    // rom_array[8578] = 32'h00006561;
    // rom_array[8579] = 32'hFFFFFFF1;
    // rom_array[8580] = 32'hFFFFFFF1;
    // rom_array[8581] = 32'h00006569;
    // rom_array[8582] = 32'h00006571;
    // rom_array[8583] = 32'hFFFFFFF1;
    // rom_array[8584] = 32'hFFFFFFF1;
    // rom_array[8585] = 32'h00006579;
    // rom_array[8586] = 32'h00006581;
    // rom_array[8587] = 32'hFFFFFFF1;
    // rom_array[8588] = 32'hFFFFFFF1;
    // rom_array[8589] = 32'h00006589;
    // rom_array[8590] = 32'h00006591;
    // rom_array[8591] = 32'h00006599;
    // rom_array[8592] = 32'h000065a1;
    // rom_array[8593] = 32'h000065a9;
    // rom_array[8594] = 32'h000065b1;
    // rom_array[8595] = 32'hFFFFFFF0;
    // rom_array[8596] = 32'hFFFFFFF0;
    // rom_array[8597] = 32'h000065b9;
    // rom_array[8598] = 32'h000065c1;
    // rom_array[8599] = 32'hFFFFFFF0;
    // rom_array[8600] = 32'hFFFFFFF0;
    // rom_array[8601] = 32'hFFFFFFF1;
    // rom_array[8602] = 32'hFFFFFFF1;
    // rom_array[8603] = 32'hFFFFFFF1;
    // rom_array[8604] = 32'hFFFFFFF1;
    // rom_array[8605] = 32'h000065c9;
    // rom_array[8606] = 32'h000065d1;
    // rom_array[8607] = 32'h000065d9;
    // rom_array[8608] = 32'h000065e1;
    // rom_array[8609] = 32'h000065e9;
    // rom_array[8610] = 32'h000065f1;
    // rom_array[8611] = 32'hFFFFFFF0;
    // rom_array[8612] = 32'hFFFFFFF0;
    // rom_array[8613] = 32'h000065f9;
    // rom_array[8614] = 32'h00006601;
    // rom_array[8615] = 32'hFFFFFFF0;
    // rom_array[8616] = 32'hFFFFFFF0;
    // rom_array[8617] = 32'h00006609;
    // rom_array[8618] = 32'h00006611;
    // rom_array[8619] = 32'h00006619;
    // rom_array[8620] = 32'h00006621;
    // rom_array[8621] = 32'h00006629;
    // rom_array[8622] = 32'h00006631;
    // rom_array[8623] = 32'h00006639;
    // rom_array[8624] = 32'h00006641;
    // rom_array[8625] = 32'h00006649;
    // rom_array[8626] = 32'h00006651;
    // rom_array[8627] = 32'h00006659;
    // rom_array[8628] = 32'h00006661;
    // rom_array[8629] = 32'h00006669;
    // rom_array[8630] = 32'h00006671;
    // rom_array[8631] = 32'h00006679;
    // rom_array[8632] = 32'h00006681;
    // rom_array[8633] = 32'h00006689;
    // rom_array[8634] = 32'h00006691;
    // rom_array[8635] = 32'h00006699;
    // rom_array[8636] = 32'h000066a1;
    // rom_array[8637] = 32'h000066a9;
    // rom_array[8638] = 32'h000066b1;
    // rom_array[8639] = 32'h000066b9;
    // rom_array[8640] = 32'h000066c1;
    // rom_array[8641] = 32'h000066c9;
    // rom_array[8642] = 32'h000066d1;
    // rom_array[8643] = 32'h000066d9;
    // rom_array[8644] = 32'h000066e1;
    // rom_array[8645] = 32'h000066e9;
    // rom_array[8646] = 32'h000066f1;
    // rom_array[8647] = 32'h000066f9;
    // rom_array[8648] = 32'h00006701;
    // rom_array[8649] = 32'h00006709;
    // rom_array[8650] = 32'h00006711;
    // rom_array[8651] = 32'h00006719;
    // rom_array[8652] = 32'h00006721;
    // rom_array[8653] = 32'h00006729;
    // rom_array[8654] = 32'h00006731;
    // rom_array[8655] = 32'h00006739;
    // rom_array[8656] = 32'h00006741;
    // rom_array[8657] = 32'h00006749;
    // rom_array[8658] = 32'h00006751;
    // rom_array[8659] = 32'hFFFFFFF0;
    // rom_array[8660] = 32'hFFFFFFF0;
    // rom_array[8661] = 32'h00006759;
    // rom_array[8662] = 32'h00006761;
    // rom_array[8663] = 32'h00006769;
    // rom_array[8664] = 32'h00006771;
    // rom_array[8665] = 32'h00006779;
    // rom_array[8666] = 32'h00006781;
    // rom_array[8667] = 32'h00006789;
    // rom_array[8668] = 32'h00006791;
    // rom_array[8669] = 32'hFFFFFFF0;
    // rom_array[8670] = 32'hFFFFFFF0;
    // rom_array[8671] = 32'hFFFFFFF0;
    // rom_array[8672] = 32'hFFFFFFF0;
    // rom_array[8673] = 32'h00006799;
    // rom_array[8674] = 32'h000067a1;
    // rom_array[8675] = 32'h000067a9;
    // rom_array[8676] = 32'h000067b1;
    // rom_array[8677] = 32'hFFFFFFF0;
    // rom_array[8678] = 32'hFFFFFFF0;
    // rom_array[8679] = 32'hFFFFFFF0;
    // rom_array[8680] = 32'hFFFFFFF0;
    // rom_array[8681] = 32'h000067b9;
    // rom_array[8682] = 32'h000067c1;
    // rom_array[8683] = 32'h000067c9;
    // rom_array[8684] = 32'h000067d1;
    // rom_array[8685] = 32'hFFFFFFF0;
    // rom_array[8686] = 32'hFFFFFFF0;
    // rom_array[8687] = 32'hFFFFFFF0;
    // rom_array[8688] = 32'hFFFFFFF0;
    // rom_array[8689] = 32'h000067d9;
    // rom_array[8690] = 32'h000067e1;
    // rom_array[8691] = 32'h000067e9;
    // rom_array[8692] = 32'h000067f1;
    // rom_array[8693] = 32'hFFFFFFF0;
    // rom_array[8694] = 32'hFFFFFFF0;
    // rom_array[8695] = 32'hFFFFFFF0;
    // rom_array[8696] = 32'hFFFFFFF0;
    // rom_array[8697] = 32'h000067f9;
    // rom_array[8698] = 32'h00006801;
    // rom_array[8699] = 32'h00006809;
    // rom_array[8700] = 32'h00006811;
    // rom_array[8701] = 32'h00006819;
    // rom_array[8702] = 32'h00006821;
    // rom_array[8703] = 32'h00006829;
    // rom_array[8704] = 32'h00006831;
    // rom_array[8705] = 32'h00006839;
    // rom_array[8706] = 32'h00006841;
    // rom_array[8707] = 32'h00006849;
    // rom_array[8708] = 32'h00006851;
    // rom_array[8709] = 32'hFFFFFFF0;
    // rom_array[8710] = 32'hFFFFFFF0;
    // rom_array[8711] = 32'hFFFFFFF0;
    // rom_array[8712] = 32'hFFFFFFF0;
    // rom_array[8713] = 32'h00006859;
    // rom_array[8714] = 32'h00006861;
    // rom_array[8715] = 32'h00006869;
    // rom_array[8716] = 32'h00006871;
    // rom_array[8717] = 32'hFFFFFFF1;
    // rom_array[8718] = 32'hFFFFFFF1;
    // rom_array[8719] = 32'h00006879;
    // rom_array[8720] = 32'h00006881;
    // rom_array[8721] = 32'hFFFFFFF1;
    // rom_array[8722] = 32'hFFFFFFF1;
    // rom_array[8723] = 32'h00006889;
    // rom_array[8724] = 32'h00006891;
    // rom_array[8725] = 32'hFFFFFFF1;
    // rom_array[8726] = 32'hFFFFFFF1;
    // rom_array[8727] = 32'h00006899;
    // rom_array[8728] = 32'h000068a1;
    // rom_array[8729] = 32'hFFFFFFF1;
    // rom_array[8730] = 32'hFFFFFFF1;
    // rom_array[8731] = 32'h000068a9;
    // rom_array[8732] = 32'h000068b1;
    // rom_array[8733] = 32'hFFFFFFF1;
    // rom_array[8734] = 32'hFFFFFFF1;
    // rom_array[8735] = 32'h000068b9;
    // rom_array[8736] = 32'h000068c1;
    // rom_array[8737] = 32'h000068c9;
    // rom_array[8738] = 32'h000068d1;
    // rom_array[8739] = 32'h000068d9;
    // rom_array[8740] = 32'h000068e1;
    // rom_array[8741] = 32'hFFFFFFF1;
    // rom_array[8742] = 32'hFFFFFFF1;
    // rom_array[8743] = 32'hFFFFFFF1;
    // rom_array[8744] = 32'hFFFFFFF1;
    // rom_array[8745] = 32'h000068e9;
    // rom_array[8746] = 32'h000068f1;
    // rom_array[8747] = 32'h000068f9;
    // rom_array[8748] = 32'h00006901;
    // rom_array[8749] = 32'hFFFFFFF1;
    // rom_array[8750] = 32'hFFFFFFF1;
    // rom_array[8751] = 32'hFFFFFFF1;
    // rom_array[8752] = 32'hFFFFFFF1;
    // rom_array[8753] = 32'h00006909;
    // rom_array[8754] = 32'h00006911;
    // rom_array[8755] = 32'h00006919;
    // rom_array[8756] = 32'h00006921;
    // rom_array[8757] = 32'hFFFFFFF0;
    // rom_array[8758] = 32'hFFFFFFF0;
    // rom_array[8759] = 32'hFFFFFFF0;
    // rom_array[8760] = 32'hFFFFFFF0;
    // rom_array[8761] = 32'h00006929;
    // rom_array[8762] = 32'h00006931;
    // rom_array[8763] = 32'h00006939;
    // rom_array[8764] = 32'h00006941;
    // rom_array[8765] = 32'hFFFFFFF0;
    // rom_array[8766] = 32'hFFFFFFF0;
    // rom_array[8767] = 32'hFFFFFFF0;
    // rom_array[8768] = 32'hFFFFFFF0;
    // rom_array[8769] = 32'h00006949;
    // rom_array[8770] = 32'h00006951;
    // rom_array[8771] = 32'h00006959;
    // rom_array[8772] = 32'h00006961;
    // rom_array[8773] = 32'hFFFFFFF1;
    // rom_array[8774] = 32'hFFFFFFF1;
    // rom_array[8775] = 32'hFFFFFFF1;
    // rom_array[8776] = 32'hFFFFFFF1;
    // rom_array[8777] = 32'h00006969;
    // rom_array[8778] = 32'h00006971;
    // rom_array[8779] = 32'h00006979;
    // rom_array[8780] = 32'h00006981;
    // rom_array[8781] = 32'hFFFFFFF1;
    // rom_array[8782] = 32'hFFFFFFF1;
    // rom_array[8783] = 32'hFFFFFFF1;
    // rom_array[8784] = 32'hFFFFFFF1;
    // rom_array[8785] = 32'h00006989;
    // rom_array[8786] = 32'h00006991;
    // rom_array[8787] = 32'h00006999;
    // rom_array[8788] = 32'h000069a1;
    // rom_array[8789] = 32'hFFFFFFF0;
    // rom_array[8790] = 32'hFFFFFFF0;
    // rom_array[8791] = 32'hFFFFFFF0;
    // rom_array[8792] = 32'hFFFFFFF0;
    // rom_array[8793] = 32'h000069a9;
    // rom_array[8794] = 32'h000069b1;
    // rom_array[8795] = 32'h000069b9;
    // rom_array[8796] = 32'h000069c1;
    // rom_array[8797] = 32'hFFFFFFF0;
    // rom_array[8798] = 32'hFFFFFFF0;
    // rom_array[8799] = 32'hFFFFFFF0;
    // rom_array[8800] = 32'hFFFFFFF0;
    // rom_array[8801] = 32'h000069c9;
    // rom_array[8802] = 32'h000069d1;
    // rom_array[8803] = 32'h000069d9;
    // rom_array[8804] = 32'h000069e1;
    // rom_array[8805] = 32'hFFFFFFF1;
    // rom_array[8806] = 32'hFFFFFFF1;
    // rom_array[8807] = 32'hFFFFFFF1;
    // rom_array[8808] = 32'hFFFFFFF1;
    // rom_array[8809] = 32'h000069e9;
    // rom_array[8810] = 32'h000069f1;
    // rom_array[8811] = 32'h000069f9;
    // rom_array[8812] = 32'h00006a01;
    // rom_array[8813] = 32'hFFFFFFF1;
    // rom_array[8814] = 32'hFFFFFFF1;
    // rom_array[8815] = 32'h00006a09;
    // rom_array[8816] = 32'h00006a11;
    // rom_array[8817] = 32'h00006a19;
    // rom_array[8818] = 32'h00006a21;
    // rom_array[8819] = 32'h00006a29;
    // rom_array[8820] = 32'h00006a31;
    // rom_array[8821] = 32'hFFFFFFF0;
    // rom_array[8822] = 32'hFFFFFFF0;
    // rom_array[8823] = 32'hFFFFFFF0;
    // rom_array[8824] = 32'hFFFFFFF0;
    // rom_array[8825] = 32'h00006a39;
    // rom_array[8826] = 32'h00006a41;
    // rom_array[8827] = 32'h00006a49;
    // rom_array[8828] = 32'h00006a51;
    // rom_array[8829] = 32'hFFFFFFF1;
    // rom_array[8830] = 32'hFFFFFFF1;
    // rom_array[8831] = 32'h00006a59;
    // rom_array[8832] = 32'h00006a61;
    // rom_array[8833] = 32'hFFFFFFF1;
    // rom_array[8834] = 32'hFFFFFFF1;
    // rom_array[8835] = 32'h00006a69;
    // rom_array[8836] = 32'h00006a71;
    // rom_array[8837] = 32'hFFFFFFF1;
    // rom_array[8838] = 32'hFFFFFFF1;
    // rom_array[8839] = 32'h00006a79;
    // rom_array[8840] = 32'h00006a81;
    // rom_array[8841] = 32'hFFFFFFF1;
    // rom_array[8842] = 32'hFFFFFFF1;
    // rom_array[8843] = 32'h00006a89;
    // rom_array[8844] = 32'h00006a91;
    // rom_array[8845] = 32'hFFFFFFF1;
    // rom_array[8846] = 32'hFFFFFFF1;
    // rom_array[8847] = 32'h00006a99;
    // rom_array[8848] = 32'h00006aa1;
    // rom_array[8849] = 32'h00006aa9;
    // rom_array[8850] = 32'h00006ab1;
    // rom_array[8851] = 32'h00006ab9;
    // rom_array[8852] = 32'h00006ac1;
    // rom_array[8853] = 32'hFFFFFFF1;
    // rom_array[8854] = 32'hFFFFFFF1;
    // rom_array[8855] = 32'hFFFFFFF1;
    // rom_array[8856] = 32'hFFFFFFF1;
    // rom_array[8857] = 32'h00006ac9;
    // rom_array[8858] = 32'h00006ad1;
    // rom_array[8859] = 32'h00006ad9;
    // rom_array[8860] = 32'h00006ae1;
    // rom_array[8861] = 32'hFFFFFFF1;
    // rom_array[8862] = 32'hFFFFFFF1;
    // rom_array[8863] = 32'hFFFFFFF1;
    // rom_array[8864] = 32'hFFFFFFF1;
    // rom_array[8865] = 32'hFFFFFFF1;
    // rom_array[8866] = 32'hFFFFFFF1;
    // rom_array[8867] = 32'hFFFFFFF1;
    // rom_array[8868] = 32'hFFFFFFF1;
    // rom_array[8869] = 32'h00006ae9;
    // rom_array[8870] = 32'h00006af1;
    // rom_array[8871] = 32'h00006af9;
    // rom_array[8872] = 32'h00006b01;
    // rom_array[8873] = 32'hFFFFFFF1;
    // rom_array[8874] = 32'hFFFFFFF1;
    // rom_array[8875] = 32'hFFFFFFF1;
    // rom_array[8876] = 32'hFFFFFFF1;
    // rom_array[8877] = 32'h00006b09;
    // rom_array[8878] = 32'h00006b11;
    // rom_array[8879] = 32'h00006b19;
    // rom_array[8880] = 32'h00006b21;
    // rom_array[8881] = 32'h00006b29;
    // rom_array[8882] = 32'h00006b31;
    // rom_array[8883] = 32'h00006b39;
    // rom_array[8884] = 32'h00006b41;
    // rom_array[8885] = 32'hFFFFFFF1;
    // rom_array[8886] = 32'hFFFFFFF1;
    // rom_array[8887] = 32'hFFFFFFF1;
    // rom_array[8888] = 32'hFFFFFFF1;
    // rom_array[8889] = 32'h00006b49;
    // rom_array[8890] = 32'h00006b51;
    // rom_array[8891] = 32'h00006b59;
    // rom_array[8892] = 32'h00006b61;
    // rom_array[8893] = 32'hFFFFFFF1;
    // rom_array[8894] = 32'hFFFFFFF1;
    // rom_array[8895] = 32'hFFFFFFF1;
    // rom_array[8896] = 32'hFFFFFFF1;
    // rom_array[8897] = 32'hFFFFFFF1;
    // rom_array[8898] = 32'hFFFFFFF1;
    // rom_array[8899] = 32'hFFFFFFF1;
    // rom_array[8900] = 32'hFFFFFFF1;
    // rom_array[8901] = 32'h00006b69;
    // rom_array[8902] = 32'h00006b71;
    // rom_array[8903] = 32'h00006b79;
    // rom_array[8904] = 32'h00006b81;
    // rom_array[8905] = 32'hFFFFFFF1;
    // rom_array[8906] = 32'hFFFFFFF1;
    // rom_array[8907] = 32'hFFFFFFF1;
    // rom_array[8908] = 32'hFFFFFFF1;
    // rom_array[8909] = 32'h00006b89;
    // rom_array[8910] = 32'h00006b91;
    // rom_array[8911] = 32'h00006b99;
    // rom_array[8912] = 32'h00006ba1;
    // rom_array[8913] = 32'h00006ba9;
    // rom_array[8914] = 32'h00006bb1;
    // rom_array[8915] = 32'h00006bb9;
    // rom_array[8916] = 32'h00006bc1;
    // rom_array[8917] = 32'hFFFFFFF0;
    // rom_array[8918] = 32'hFFFFFFF0;
    // rom_array[8919] = 32'hFFFFFFF0;
    // rom_array[8920] = 32'hFFFFFFF0;
    // rom_array[8921] = 32'h00006bc9;
    // rom_array[8922] = 32'h00006bd1;
    // rom_array[8923] = 32'h00006bd9;
    // rom_array[8924] = 32'h00006be1;
    // rom_array[8925] = 32'hFFFFFFF0;
    // rom_array[8926] = 32'hFFFFFFF0;
    // rom_array[8927] = 32'hFFFFFFF0;
    // rom_array[8928] = 32'hFFFFFFF0;
    // rom_array[8929] = 32'h00006be9;
    // rom_array[8930] = 32'h00006bf1;
    // rom_array[8931] = 32'h00006bf9;
    // rom_array[8932] = 32'h00006c01;
    // rom_array[8933] = 32'hFFFFFFF0;
    // rom_array[8934] = 32'hFFFFFFF0;
    // rom_array[8935] = 32'hFFFFFFF0;
    // rom_array[8936] = 32'hFFFFFFF0;
    // rom_array[8937] = 32'h00006c09;
    // rom_array[8938] = 32'h00006c11;
    // rom_array[8939] = 32'h00006c19;
    // rom_array[8940] = 32'h00006c21;
    // rom_array[8941] = 32'hFFFFFFF0;
    // rom_array[8942] = 32'hFFFFFFF0;
    // rom_array[8943] = 32'hFFFFFFF0;
    // rom_array[8944] = 32'hFFFFFFF0;
    // rom_array[8945] = 32'h00006c29;
    // rom_array[8946] = 32'h00006c31;
    // rom_array[8947] = 32'h00006c39;
    // rom_array[8948] = 32'h00006c41;
    // rom_array[8949] = 32'hFFFFFFF1;
    // rom_array[8950] = 32'hFFFFFFF1;
    // rom_array[8951] = 32'hFFFFFFF1;
    // rom_array[8952] = 32'hFFFFFFF1;
    // rom_array[8953] = 32'h00006c49;
    // rom_array[8954] = 32'h00006c51;
    // rom_array[8955] = 32'h00006c59;
    // rom_array[8956] = 32'h00006c61;
    // rom_array[8957] = 32'h00006c69;
    // rom_array[8958] = 32'h00006c71;
    // rom_array[8959] = 32'h00006c79;
    // rom_array[8960] = 32'h00006c81;
    // rom_array[8961] = 32'hFFFFFFF1;
    // rom_array[8962] = 32'hFFFFFFF1;
    // rom_array[8963] = 32'hFFFFFFF1;
    // rom_array[8964] = 32'hFFFFFFF1;
    // rom_array[8965] = 32'h00006c89;
    // rom_array[8966] = 32'h00006c91;
    // rom_array[8967] = 32'h00006c99;
    // rom_array[8968] = 32'h00006ca1;
    // rom_array[8969] = 32'h00006ca9;
    // rom_array[8970] = 32'h00006cb1;
    // rom_array[8971] = 32'h00006cb9;
    // rom_array[8972] = 32'h00006cc1;
    // rom_array[8973] = 32'h00006cc9;
    // rom_array[8974] = 32'h00006cd1;
    // rom_array[8975] = 32'h00006cd9;
    // rom_array[8976] = 32'h00006ce1;
    // rom_array[8977] = 32'h00006ce9;
    // rom_array[8978] = 32'h00006cf1;
    // rom_array[8979] = 32'h00006cf9;
    // rom_array[8980] = 32'h00006d01;
    // rom_array[8981] = 32'hFFFFFFF0;
    // rom_array[8982] = 32'hFFFFFFF0;
    // rom_array[8983] = 32'hFFFFFFF0;
    // rom_array[8984] = 32'hFFFFFFF0;
    // rom_array[8985] = 32'h00006d09;
    // rom_array[8986] = 32'h00006d11;
    // rom_array[8987] = 32'hFFFFFFF0;
    // rom_array[8988] = 32'hFFFFFFF0;
    // rom_array[8989] = 32'hFFFFFFF0;
    // rom_array[8990] = 32'hFFFFFFF0;
    // rom_array[8991] = 32'hFFFFFFF0;
    // rom_array[8992] = 32'hFFFFFFF0;
    // rom_array[8993] = 32'h00006d19;
    // rom_array[8994] = 32'h00006d21;
    // rom_array[8995] = 32'h00006d29;
    // rom_array[8996] = 32'h00006d31;
    // rom_array[8997] = 32'hFFFFFFF1;
    // rom_array[8998] = 32'hFFFFFFF1;
    // rom_array[8999] = 32'hFFFFFFF1;
    // rom_array[9000] = 32'hFFFFFFF1;
    // rom_array[9001] = 32'h00006d39;
    // rom_array[9002] = 32'h00006d41;
    // rom_array[9003] = 32'h00006d49;
    // rom_array[9004] = 32'h00006d51;
    // rom_array[9005] = 32'hFFFFFFF1;
    // rom_array[9006] = 32'hFFFFFFF1;
    // rom_array[9007] = 32'hFFFFFFF1;
    // rom_array[9008] = 32'hFFFFFFF1;
    // rom_array[9009] = 32'h00006d59;
    // rom_array[9010] = 32'h00006d61;
    // rom_array[9011] = 32'h00006d69;
    // rom_array[9012] = 32'h00006d71;
    // rom_array[9013] = 32'hFFFFFFF1;
    // rom_array[9014] = 32'hFFFFFFF1;
    // rom_array[9015] = 32'hFFFFFFF1;
    // rom_array[9016] = 32'hFFFFFFF1;
    // rom_array[9017] = 32'h00006d79;
    // rom_array[9018] = 32'h00006d81;
    // rom_array[9019] = 32'h00006d89;
    // rom_array[9020] = 32'h00006d91;
    // rom_array[9021] = 32'hFFFFFFF1;
    // rom_array[9022] = 32'hFFFFFFF1;
    // rom_array[9023] = 32'hFFFFFFF1;
    // rom_array[9024] = 32'hFFFFFFF1;
    // rom_array[9025] = 32'h00006d99;
    // rom_array[9026] = 32'h00006da1;
    // rom_array[9027] = 32'h00006da9;
    // rom_array[9028] = 32'h00006db1;
    // rom_array[9029] = 32'h00006db9;
    // rom_array[9030] = 32'h00006dc1;
    // rom_array[9031] = 32'hFFFFFFF0;
    // rom_array[9032] = 32'hFFFFFFF0;
    // rom_array[9033] = 32'h00006dc9;
    // rom_array[9034] = 32'h00006dd1;
    // rom_array[9035] = 32'h00006dd9;
    // rom_array[9036] = 32'h00006de1;
    // rom_array[9037] = 32'hFFFFFFF0;
    // rom_array[9038] = 32'hFFFFFFF0;
    // rom_array[9039] = 32'hFFFFFFF0;
    // rom_array[9040] = 32'hFFFFFFF0;
    // rom_array[9041] = 32'h00006de9;
    // rom_array[9042] = 32'h00006df1;
    // rom_array[9043] = 32'hFFFFFFF0;
    // rom_array[9044] = 32'hFFFFFFF0;
    // rom_array[9045] = 32'h00006df9;
    // rom_array[9046] = 32'h00006e01;
    // rom_array[9047] = 32'hFFFFFFF0;
    // rom_array[9048] = 32'hFFFFFFF0;
    // rom_array[9049] = 32'h00006e09;
    // rom_array[9050] = 32'h00006e11;
    // rom_array[9051] = 32'h00006e19;
    // rom_array[9052] = 32'h00006e21;
    // rom_array[9053] = 32'hFFFFFFF0;
    // rom_array[9054] = 32'hFFFFFFF0;
    // rom_array[9055] = 32'hFFFFFFF0;
    // rom_array[9056] = 32'hFFFFFFF0;
    // rom_array[9057] = 32'h00006e29;
    // rom_array[9058] = 32'h00006e31;
    // rom_array[9059] = 32'h00006e39;
    // rom_array[9060] = 32'h00006e41;
    // rom_array[9061] = 32'h00006e49;
    // rom_array[9062] = 32'h00006e51;
    // rom_array[9063] = 32'hFFFFFFF1;
    // rom_array[9064] = 32'hFFFFFFF1;
    // rom_array[9065] = 32'h00006e59;
    // rom_array[9066] = 32'h00006e61;
    // rom_array[9067] = 32'hFFFFFFF1;
    // rom_array[9068] = 32'hFFFFFFF1;
    // rom_array[9069] = 32'h00006e69;
    // rom_array[9070] = 32'h00006e71;
    // rom_array[9071] = 32'hFFFFFFF1;
    // rom_array[9072] = 32'hFFFFFFF1;
    // rom_array[9073] = 32'h00006e79;
    // rom_array[9074] = 32'h00006e81;
    // rom_array[9075] = 32'h00006e89;
    // rom_array[9076] = 32'h00006e91;
    // rom_array[9077] = 32'hFFFFFFF1;
    // rom_array[9078] = 32'hFFFFFFF1;
    // rom_array[9079] = 32'hFFFFFFF1;
    // rom_array[9080] = 32'hFFFFFFF1;
    // rom_array[9081] = 32'h00006e99;
    // rom_array[9082] = 32'h00006ea1;
    // rom_array[9083] = 32'hFFFFFFF0;
    // rom_array[9084] = 32'hFFFFFFF0;
    // rom_array[9085] = 32'h00006ea9;
    // rom_array[9086] = 32'h00006eb1;
    // rom_array[9087] = 32'hFFFFFFF0;
    // rom_array[9088] = 32'hFFFFFFF0;
    // rom_array[9089] = 32'h00006eb9;
    // rom_array[9090] = 32'h00006ec1;
    // rom_array[9091] = 32'hFFFFFFF0;
    // rom_array[9092] = 32'hFFFFFFF0;
    // rom_array[9093] = 32'h00006ec9;
    // rom_array[9094] = 32'h00006ed1;
    // rom_array[9095] = 32'hFFFFFFF0;
    // rom_array[9096] = 32'hFFFFFFF0;
    // rom_array[9097] = 32'h00006ed9;
    // rom_array[9098] = 32'h00006ee1;
    // rom_array[9099] = 32'h00006ee9;
    // rom_array[9100] = 32'h00006ef1;
    // rom_array[9101] = 32'hFFFFFFF1;
    // rom_array[9102] = 32'hFFFFFFF1;
    // rom_array[9103] = 32'hFFFFFFF1;
    // rom_array[9104] = 32'hFFFFFFF1;
    // rom_array[9105] = 32'h00006ef9;
    // rom_array[9106] = 32'h00006f01;
    // rom_array[9107] = 32'hFFFFFFF0;
    // rom_array[9108] = 32'hFFFFFFF0;
    // rom_array[9109] = 32'h00006f09;
    // rom_array[9110] = 32'h00006f11;
    // rom_array[9111] = 32'hFFFFFFF0;
    // rom_array[9112] = 32'hFFFFFFF0;
    // rom_array[9113] = 32'h00006f19;
    // rom_array[9114] = 32'h00006f21;
    // rom_array[9115] = 32'hFFFFFFF0;
    // rom_array[9116] = 32'hFFFFFFF0;
    // rom_array[9117] = 32'h00006f29;
    // rom_array[9118] = 32'h00006f31;
    // rom_array[9119] = 32'hFFFFFFF0;
    // rom_array[9120] = 32'hFFFFFFF0;
    // rom_array[9121] = 32'h00006f39;
    // rom_array[9122] = 32'h00006f41;
    // rom_array[9123] = 32'hFFFFFFF0;
    // rom_array[9124] = 32'hFFFFFFF0;
    // rom_array[9125] = 32'h00006f49;
    // rom_array[9126] = 32'h00006f51;
    // rom_array[9127] = 32'hFFFFFFF0;
    // rom_array[9128] = 32'hFFFFFFF0;
    // rom_array[9129] = 32'h00006f59;
    // rom_array[9130] = 32'h00006f61;
    // rom_array[9131] = 32'hFFFFFFF0;
    // rom_array[9132] = 32'hFFFFFFF0;
    // rom_array[9133] = 32'h00006f69;
    // rom_array[9134] = 32'h00006f71;
    // rom_array[9135] = 32'h00006f79;
    // rom_array[9136] = 32'h00006f81;
    // rom_array[9137] = 32'hFFFFFFF0;
    // rom_array[9138] = 32'hFFFFFFF0;
    // rom_array[9139] = 32'hFFFFFFF0;
    // rom_array[9140] = 32'hFFFFFFF0;
    // rom_array[9141] = 32'h00006f89;
    // rom_array[9142] = 32'h00006f91;
    // rom_array[9143] = 32'h00006f99;
    // rom_array[9144] = 32'h00006fa1;
    // rom_array[9145] = 32'h00006fa9;
    // rom_array[9146] = 32'h00006fb1;
    // rom_array[9147] = 32'hFFFFFFF1;
    // rom_array[9148] = 32'hFFFFFFF1;
    // rom_array[9149] = 32'h00006fb9;
    // rom_array[9150] = 32'h00006fc1;
    // rom_array[9151] = 32'hFFFFFFF1;
    // rom_array[9152] = 32'hFFFFFFF1;
    // rom_array[9153] = 32'hFFFFFFF0;
    // rom_array[9154] = 32'hFFFFFFF0;
    // rom_array[9155] = 32'hFFFFFFF0;
    // rom_array[9156] = 32'hFFFFFFF0;
    // rom_array[9157] = 32'h00006fc9;
    // rom_array[9158] = 32'h00006fd1;
    // rom_array[9159] = 32'h00006fd9;
    // rom_array[9160] = 32'h00006fe1;
    // rom_array[9161] = 32'h00006fe9;
    // rom_array[9162] = 32'h00006ff1;
    // rom_array[9163] = 32'hFFFFFFF1;
    // rom_array[9164] = 32'hFFFFFFF1;
    // rom_array[9165] = 32'h00006ff9;
    // rom_array[9166] = 32'h00007001;
    // rom_array[9167] = 32'h00007009;
    // rom_array[9168] = 32'h00007011;
    // rom_array[9169] = 32'h00007019;
    // rom_array[9170] = 32'h00007021;
    // rom_array[9171] = 32'hFFFFFFF0;
    // rom_array[9172] = 32'hFFFFFFF0;
    // rom_array[9173] = 32'hFFFFFFF0;
    // rom_array[9174] = 32'hFFFFFFF0;
    // rom_array[9175] = 32'hFFFFFFF0;
    // rom_array[9176] = 32'hFFFFFFF0;
    // rom_array[9177] = 32'hFFFFFFF1;
    // rom_array[9178] = 32'hFFFFFFF1;
    // rom_array[9179] = 32'hFFFFFFF1;
    // rom_array[9180] = 32'hFFFFFFF1;
    // rom_array[9181] = 32'h00007029;
    // rom_array[9182] = 32'h00007031;
    // rom_array[9183] = 32'h00007039;
    // rom_array[9184] = 32'h00007041;
    // rom_array[9185] = 32'hFFFFFFF1;
    // rom_array[9186] = 32'hFFFFFFF1;
    // rom_array[9187] = 32'hFFFFFFF1;
    // rom_array[9188] = 32'hFFFFFFF1;
    // rom_array[9189] = 32'h00007049;
    // rom_array[9190] = 32'h00007051;
    // rom_array[9191] = 32'h00007059;
    // rom_array[9192] = 32'h00007061;
    // rom_array[9193] = 32'h00007069;
    // rom_array[9194] = 32'h00007071;
    // rom_array[9195] = 32'h00007079;
    // rom_array[9196] = 32'h00007081;
    // rom_array[9197] = 32'hFFFFFFF1;
    // rom_array[9198] = 32'hFFFFFFF1;
    // rom_array[9199] = 32'h00007089;
    // rom_array[9200] = 32'h00007091;
    // rom_array[9201] = 32'hFFFFFFF1;
    // rom_array[9202] = 32'hFFFFFFF1;
    // rom_array[9203] = 32'hFFFFFFF1;
    // rom_array[9204] = 32'hFFFFFFF1;
    // rom_array[9205] = 32'h00007099;
    // rom_array[9206] = 32'h000070a1;
    // rom_array[9207] = 32'h000070a9;
    // rom_array[9208] = 32'h000070b1;
    // rom_array[9209] = 32'hFFFFFFF1;
    // rom_array[9210] = 32'hFFFFFFF1;
    // rom_array[9211] = 32'h000070b9;
    // rom_array[9212] = 32'h000070c1;
    // rom_array[9213] = 32'h000070c9;
    // rom_array[9214] = 32'h000070d1;
    // rom_array[9215] = 32'h000070d9;
    // rom_array[9216] = 32'h000070e1;
    // rom_array[9217] = 32'h000070e9;
    // rom_array[9218] = 32'h000070f1;
    // rom_array[9219] = 32'hFFFFFFF0;
    // rom_array[9220] = 32'hFFFFFFF0;
    // rom_array[9221] = 32'h000070f9;
    // rom_array[9222] = 32'h00007101;
    // rom_array[9223] = 32'hFFFFFFF0;
    // rom_array[9224] = 32'hFFFFFFF0;
    // rom_array[9225] = 32'h00007109;
    // rom_array[9226] = 32'h00007111;
    // rom_array[9227] = 32'hFFFFFFF0;
    // rom_array[9228] = 32'hFFFFFFF0;
    // rom_array[9229] = 32'h00007119;
    // rom_array[9230] = 32'h00007121;
    // rom_array[9231] = 32'hFFFFFFF0;
    // rom_array[9232] = 32'hFFFFFFF0;
    // rom_array[9233] = 32'h00007129;
    // rom_array[9234] = 32'h00007131;
    // rom_array[9235] = 32'h00007139;
    // rom_array[9236] = 32'h00007141;
    // rom_array[9237] = 32'hFFFFFFF0;
    // rom_array[9238] = 32'hFFFFFFF0;
    // rom_array[9239] = 32'hFFFFFFF0;
    // rom_array[9240] = 32'hFFFFFFF0;
    // rom_array[9241] = 32'h00007149;
    // rom_array[9242] = 32'h00007151;
    // rom_array[9243] = 32'hFFFFFFF0;
    // rom_array[9244] = 32'hFFFFFFF0;
    // rom_array[9245] = 32'hFFFFFFF0;
    // rom_array[9246] = 32'hFFFFFFF0;
    // rom_array[9247] = 32'hFFFFFFF0;
    // rom_array[9248] = 32'hFFFFFFF0;
    // rom_array[9249] = 32'h00007159;
    // rom_array[9250] = 32'h00007161;
    // rom_array[9251] = 32'h00007169;
    // rom_array[9252] = 32'h00007171;
    // rom_array[9253] = 32'hFFFFFFF1;
    // rom_array[9254] = 32'hFFFFFFF1;
    // rom_array[9255] = 32'hFFFFFFF1;
    // rom_array[9256] = 32'hFFFFFFF1;
    // rom_array[9257] = 32'h00007179;
    // rom_array[9258] = 32'h00007181;
    // rom_array[9259] = 32'h00007189;
    // rom_array[9260] = 32'h00007191;
    // rom_array[9261] = 32'hFFFFFFF1;
    // rom_array[9262] = 32'hFFFFFFF1;
    // rom_array[9263] = 32'hFFFFFFF1;
    // rom_array[9264] = 32'hFFFFFFF1;
    // rom_array[9265] = 32'h00007199;
    // rom_array[9266] = 32'h000071a1;
    // rom_array[9267] = 32'h000071a9;
    // rom_array[9268] = 32'h000071b1;
    // rom_array[9269] = 32'hFFFFFFF1;
    // rom_array[9270] = 32'hFFFFFFF1;
    // rom_array[9271] = 32'hFFFFFFF1;
    // rom_array[9272] = 32'hFFFFFFF1;
    // rom_array[9273] = 32'h000071b9;
    // rom_array[9274] = 32'h000071c1;
    // rom_array[9275] = 32'h000071c9;
    // rom_array[9276] = 32'h000071d1;
    // rom_array[9277] = 32'hFFFFFFF1;
    // rom_array[9278] = 32'hFFFFFFF1;
    // rom_array[9279] = 32'hFFFFFFF1;
    // rom_array[9280] = 32'hFFFFFFF1;
    // rom_array[9281] = 32'h000071d9;
    // rom_array[9282] = 32'h000071e1;
    // rom_array[9283] = 32'h000071e9;
    // rom_array[9284] = 32'h000071f1;
    // rom_array[9285] = 32'hFFFFFFF1;
    // rom_array[9286] = 32'hFFFFFFF1;
    // rom_array[9287] = 32'h000071f9;
    // rom_array[9288] = 32'h00007201;
    // rom_array[9289] = 32'h00007209;
    // rom_array[9290] = 32'h00007211;
    // rom_array[9291] = 32'h00007219;
    // rom_array[9292] = 32'h00007221;
    // rom_array[9293] = 32'hFFFFFFF0;
    // rom_array[9294] = 32'hFFFFFFF0;
    // rom_array[9295] = 32'hFFFFFFF0;
    // rom_array[9296] = 32'hFFFFFFF0;
    // rom_array[9297] = 32'h00007229;
    // rom_array[9298] = 32'h00007231;
    // rom_array[9299] = 32'h00007239;
    // rom_array[9300] = 32'h00007241;
    // rom_array[9301] = 32'hFFFFFFF0;
    // rom_array[9302] = 32'hFFFFFFF0;
    // rom_array[9303] = 32'hFFFFFFF0;
    // rom_array[9304] = 32'hFFFFFFF0;
    // rom_array[9305] = 32'h00007249;
    // rom_array[9306] = 32'h00007251;
    // rom_array[9307] = 32'h00007259;
    // rom_array[9308] = 32'h00007261;
    // rom_array[9309] = 32'h00007269;
    // rom_array[9310] = 32'h00007271;
    // rom_array[9311] = 32'hFFFFFFF1;
    // rom_array[9312] = 32'hFFFFFFF1;
    // rom_array[9313] = 32'h00007279;
    // rom_array[9314] = 32'h00007281;
    // rom_array[9315] = 32'h00007289;
    // rom_array[9316] = 32'h00007291;
    // rom_array[9317] = 32'hFFFFFFF1;
    // rom_array[9318] = 32'hFFFFFFF1;
    // rom_array[9319] = 32'hFFFFFFF1;
    // rom_array[9320] = 32'hFFFFFFF1;
    // rom_array[9321] = 32'h00007299;
    // rom_array[9322] = 32'h000072a1;
    // rom_array[9323] = 32'hFFFFFFF0;
    // rom_array[9324] = 32'hFFFFFFF0;
    // rom_array[9325] = 32'h000072a9;
    // rom_array[9326] = 32'h000072b1;
    // rom_array[9327] = 32'hFFFFFFF0;
    // rom_array[9328] = 32'hFFFFFFF0;
    // rom_array[9329] = 32'h000072b9;
    // rom_array[9330] = 32'h000072c1;
    // rom_array[9331] = 32'hFFFFFFF0;
    // rom_array[9332] = 32'hFFFFFFF0;
    // rom_array[9333] = 32'h000072c9;
    // rom_array[9334] = 32'h000072d1;
    // rom_array[9335] = 32'hFFFFFFF0;
    // rom_array[9336] = 32'hFFFFFFF0;
    // rom_array[9337] = 32'h000072d9;
    // rom_array[9338] = 32'h000072e1;
    // rom_array[9339] = 32'h000072e9;
    // rom_array[9340] = 32'h000072f1;
    // rom_array[9341] = 32'hFFFFFFF1;
    // rom_array[9342] = 32'hFFFFFFF1;
    // rom_array[9343] = 32'hFFFFFFF1;
    // rom_array[9344] = 32'hFFFFFFF1;
    // rom_array[9345] = 32'h000072f9;
    // rom_array[9346] = 32'h00007301;
    // rom_array[9347] = 32'hFFFFFFF0;
    // rom_array[9348] = 32'hFFFFFFF0;
    // rom_array[9349] = 32'h00007309;
    // rom_array[9350] = 32'h00007311;
    // rom_array[9351] = 32'hFFFFFFF0;
    // rom_array[9352] = 32'hFFFFFFF0;
    // rom_array[9353] = 32'hFFFFFFF1;
    // rom_array[9354] = 32'hFFFFFFF1;
    // rom_array[9355] = 32'h00007319;
    // rom_array[9356] = 32'h00007321;
    // rom_array[9357] = 32'hFFFFFFF1;
    // rom_array[9358] = 32'hFFFFFFF1;
    // rom_array[9359] = 32'h00007329;
    // rom_array[9360] = 32'h00007331;
    // rom_array[9361] = 32'hFFFFFFF1;
    // rom_array[9362] = 32'hFFFFFFF1;
    // rom_array[9363] = 32'h00007339;
    // rom_array[9364] = 32'h00007341;
    // rom_array[9365] = 32'hFFFFFFF1;
    // rom_array[9366] = 32'hFFFFFFF1;
    // rom_array[9367] = 32'h00007349;
    // rom_array[9368] = 32'h00007351;
    // rom_array[9369] = 32'h00007359;
    // rom_array[9370] = 32'h00007361;
    // rom_array[9371] = 32'hFFFFFFF1;
    // rom_array[9372] = 32'hFFFFFFF1;
    // rom_array[9373] = 32'h00007369;
    // rom_array[9374] = 32'h00007371;
    // rom_array[9375] = 32'hFFFFFFF1;
    // rom_array[9376] = 32'hFFFFFFF1;
    // rom_array[9377] = 32'h00007379;
    // rom_array[9378] = 32'h00007381;
    // rom_array[9379] = 32'hFFFFFFF1;
    // rom_array[9380] = 32'hFFFFFFF1;
    // rom_array[9381] = 32'h00007389;
    // rom_array[9382] = 32'h00007391;
    // rom_array[9383] = 32'hFFFFFFF1;
    // rom_array[9384] = 32'hFFFFFFF1;
    // rom_array[9385] = 32'hFFFFFFF1;
    // rom_array[9386] = 32'hFFFFFFF1;
    // rom_array[9387] = 32'h00007399;
    // rom_array[9388] = 32'h000073a1;
    // rom_array[9389] = 32'hFFFFFFF1;
    // rom_array[9390] = 32'hFFFFFFF1;
    // rom_array[9391] = 32'h000073a9;
    // rom_array[9392] = 32'h000073b1;
    // rom_array[9393] = 32'hFFFFFFF1;
    // rom_array[9394] = 32'hFFFFFFF1;
    // rom_array[9395] = 32'h000073b9;
    // rom_array[9396] = 32'h000073c1;
    // rom_array[9397] = 32'hFFFFFFF1;
    // rom_array[9398] = 32'hFFFFFFF1;
    // rom_array[9399] = 32'h000073c9;
    // rom_array[9400] = 32'h000073d1;
    // rom_array[9401] = 32'h000073d9;
    // rom_array[9402] = 32'h000073e1;
    // rom_array[9403] = 32'hFFFFFFF1;
    // rom_array[9404] = 32'hFFFFFFF1;
    // rom_array[9405] = 32'h000073e9;
    // rom_array[9406] = 32'h000073f1;
    // rom_array[9407] = 32'hFFFFFFF1;
    // rom_array[9408] = 32'hFFFFFFF1;
    // rom_array[9409] = 32'h000073f9;
    // rom_array[9410] = 32'h00007401;
    // rom_array[9411] = 32'hFFFFFFF1;
    // rom_array[9412] = 32'hFFFFFFF1;
    // rom_array[9413] = 32'h00007409;
    // rom_array[9414] = 32'h00007411;
    // rom_array[9415] = 32'hFFFFFFF1;
    // rom_array[9416] = 32'hFFFFFFF1;
    // rom_array[9417] = 32'h00007419;
    // rom_array[9418] = 32'h00007421;
    // rom_array[9419] = 32'hFFFFFFF0;
    // rom_array[9420] = 32'hFFFFFFF0;
    // rom_array[9421] = 32'h00007429;
    // rom_array[9422] = 32'h00007431;
    // rom_array[9423] = 32'hFFFFFFF0;
    // rom_array[9424] = 32'hFFFFFFF0;
    // rom_array[9425] = 32'h00007439;
    // rom_array[9426] = 32'h00007441;
    // rom_array[9427] = 32'hFFFFFFF0;
    // rom_array[9428] = 32'hFFFFFFF0;
    // rom_array[9429] = 32'h00007449;
    // rom_array[9430] = 32'h00007451;
    // rom_array[9431] = 32'hFFFFFFF0;
    // rom_array[9432] = 32'hFFFFFFF0;
    // rom_array[9433] = 32'h00007459;
    // rom_array[9434] = 32'h00007461;
    // rom_array[9435] = 32'hFFFFFFF0;
    // rom_array[9436] = 32'hFFFFFFF0;
    // rom_array[9437] = 32'h00007469;
    // rom_array[9438] = 32'h00007471;
    // rom_array[9439] = 32'hFFFFFFF0;
    // rom_array[9440] = 32'hFFFFFFF0;
    // rom_array[9441] = 32'h00007479;
    // rom_array[9442] = 32'h00007481;
    // rom_array[9443] = 32'hFFFFFFF0;
    // rom_array[9444] = 32'hFFFFFFF0;
    // rom_array[9445] = 32'h00007489;
    // rom_array[9446] = 32'h00007491;
    // rom_array[9447] = 32'hFFFFFFF0;
    // rom_array[9448] = 32'hFFFFFFF0;
    // rom_array[9449] = 32'h00007499;
    // rom_array[9450] = 32'h000074a1;
    // rom_array[9451] = 32'h000074a9;
    // rom_array[9452] = 32'h000074b1;
    // rom_array[9453] = 32'hFFFFFFF0;
    // rom_array[9454] = 32'hFFFFFFF0;
    // rom_array[9455] = 32'hFFFFFFF0;
    // rom_array[9456] = 32'hFFFFFFF0;
    // rom_array[9457] = 32'h000074b9;
    // rom_array[9458] = 32'h000074c1;
    // rom_array[9459] = 32'h000074c9;
    // rom_array[9460] = 32'h000074d1;
    // rom_array[9461] = 32'hFFFFFFF0;
    // rom_array[9462] = 32'hFFFFFFF0;
    // rom_array[9463] = 32'hFFFFFFF0;
    // rom_array[9464] = 32'hFFFFFFF0;
    // rom_array[9465] = 32'h000074d9;
    // rom_array[9466] = 32'h000074e1;
    // rom_array[9467] = 32'hFFFFFFF0;
    // rom_array[9468] = 32'hFFFFFFF0;
    // rom_array[9469] = 32'hFFFFFFF0;
    // rom_array[9470] = 32'hFFFFFFF0;
    // rom_array[9471] = 32'hFFFFFFF0;
    // rom_array[9472] = 32'hFFFFFFF0;
    // rom_array[9473] = 32'hFFFFFFF0;
    // rom_array[9474] = 32'hFFFFFFF0;
    // rom_array[9475] = 32'h000074e9;
    // rom_array[9476] = 32'h000074f1;
    // rom_array[9477] = 32'hFFFFFFF0;
    // rom_array[9478] = 32'hFFFFFFF0;
    // rom_array[9479] = 32'hFFFFFFF0;
    // rom_array[9480] = 32'hFFFFFFF0;
    // rom_array[9481] = 32'h000074f9;
    // rom_array[9482] = 32'h00007501;
    // rom_array[9483] = 32'h00007509;
    // rom_array[9484] = 32'h00007511;
    // rom_array[9485] = 32'hFFFFFFF0;
    // rom_array[9486] = 32'hFFFFFFF0;
    // rom_array[9487] = 32'hFFFFFFF0;
    // rom_array[9488] = 32'hFFFFFFF0;
    // rom_array[9489] = 32'h00007519;
    // rom_array[9490] = 32'h00007521;
    // rom_array[9491] = 32'h00007529;
    // rom_array[9492] = 32'h00007531;
    // rom_array[9493] = 32'h00007539;
    // rom_array[9494] = 32'h00007541;
    // rom_array[9495] = 32'hFFFFFFF1;
    // rom_array[9496] = 32'hFFFFFFF1;
    // rom_array[9497] = 32'h00007549;
    // rom_array[9498] = 32'h00007551;
    // rom_array[9499] = 32'h00007559;
    // rom_array[9500] = 32'h00007561;
    // rom_array[9501] = 32'hFFFFFFF1;
    // rom_array[9502] = 32'hFFFFFFF1;
    // rom_array[9503] = 32'hFFFFFFF1;
    // rom_array[9504] = 32'hFFFFFFF1;
    // rom_array[9505] = 32'h00007569;
    // rom_array[9506] = 32'h00007571;
    // rom_array[9507] = 32'hFFFFFFF1;
    // rom_array[9508] = 32'hFFFFFFF1;
    // rom_array[9509] = 32'h00007579;
    // rom_array[9510] = 32'h00007581;
    // rom_array[9511] = 32'hFFFFFFF1;
    // rom_array[9512] = 32'hFFFFFFF1;
    // rom_array[9513] = 32'h00007589;
    // rom_array[9514] = 32'h00007591;
    // rom_array[9515] = 32'h00007599;
    // rom_array[9516] = 32'h000075a1;
    // rom_array[9517] = 32'hFFFFFFF0;
    // rom_array[9518] = 32'hFFFFFFF0;
    // rom_array[9519] = 32'hFFFFFFF0;
    // rom_array[9520] = 32'hFFFFFFF0;
    // rom_array[9521] = 32'h000075a9;
    // rom_array[9522] = 32'h000075b1;
    // rom_array[9523] = 32'h000075b9;
    // rom_array[9524] = 32'h000075c1;
    // rom_array[9525] = 32'hFFFFFFF0;
    // rom_array[9526] = 32'hFFFFFFF0;
    // rom_array[9527] = 32'hFFFFFFF0;
    // rom_array[9528] = 32'hFFFFFFF0;
    // rom_array[9529] = 32'h000075c9;
    // rom_array[9530] = 32'h000075d1;
    // rom_array[9531] = 32'h000075d9;
    // rom_array[9532] = 32'h000075e1;
    // rom_array[9533] = 32'hFFFFFFF1;
    // rom_array[9534] = 32'hFFFFFFF1;
    // rom_array[9535] = 32'hFFFFFFF1;
    // rom_array[9536] = 32'hFFFFFFF1;
    // rom_array[9537] = 32'h000075e9;
    // rom_array[9538] = 32'h000075f1;
    // rom_array[9539] = 32'h000075f9;
    // rom_array[9540] = 32'h00007601;
    // rom_array[9541] = 32'hFFFFFFF1;
    // rom_array[9542] = 32'hFFFFFFF1;
    // rom_array[9543] = 32'hFFFFFFF1;
    // rom_array[9544] = 32'hFFFFFFF1;
    // rom_array[9545] = 32'h00007609;
    // rom_array[9546] = 32'h00007611;
    // rom_array[9547] = 32'h00007619;
    // rom_array[9548] = 32'h00007621;
    // rom_array[9549] = 32'hFFFFFFF1;
    // rom_array[9550] = 32'hFFFFFFF1;
    // rom_array[9551] = 32'hFFFFFFF1;
    // rom_array[9552] = 32'hFFFFFFF1;
    // rom_array[9553] = 32'h00007629;
    // rom_array[9554] = 32'h00007631;
    // rom_array[9555] = 32'h00007639;
    // rom_array[9556] = 32'h00007641;
    // rom_array[9557] = 32'hFFFFFFF1;
    // rom_array[9558] = 32'hFFFFFFF1;
    // rom_array[9559] = 32'hFFFFFFF1;
    // rom_array[9560] = 32'hFFFFFFF1;
    // rom_array[9561] = 32'h00007649;
    // rom_array[9562] = 32'h00007651;
    // rom_array[9563] = 32'h00007659;
    // rom_array[9564] = 32'h00007661;
    // rom_array[9565] = 32'hFFFFFFF0;
    // rom_array[9566] = 32'hFFFFFFF0;
    // rom_array[9567] = 32'hFFFFFFF0;
    // rom_array[9568] = 32'hFFFFFFF0;
    // rom_array[9569] = 32'h00007669;
    // rom_array[9570] = 32'h00007671;
    // rom_array[9571] = 32'h00007679;
    // rom_array[9572] = 32'h00007681;
    // rom_array[9573] = 32'hFFFFFFF0;
    // rom_array[9574] = 32'hFFFFFFF0;
    // rom_array[9575] = 32'hFFFFFFF0;
    // rom_array[9576] = 32'hFFFFFFF0;
    // rom_array[9577] = 32'h00007689;
    // rom_array[9578] = 32'h00007691;
    // rom_array[9579] = 32'h00007699;
    // rom_array[9580] = 32'h000076a1;
    // rom_array[9581] = 32'h000076a9;
    // rom_array[9582] = 32'h000076b1;
    // rom_array[9583] = 32'hFFFFFFF1;
    // rom_array[9584] = 32'hFFFFFFF1;
    // rom_array[9585] = 32'h000076b9;
    // rom_array[9586] = 32'h000076c1;
    // rom_array[9587] = 32'h000076c9;
    // rom_array[9588] = 32'h000076d1;
    // rom_array[9589] = 32'hFFFFFFF1;
    // rom_array[9590] = 32'hFFFFFFF1;
    // rom_array[9591] = 32'hFFFFFFF1;
    // rom_array[9592] = 32'hFFFFFFF1;
    // rom_array[9593] = 32'h000076d9;
    // rom_array[9594] = 32'h000076e1;
    // rom_array[9595] = 32'h000076e9;
    // rom_array[9596] = 32'h000076f1;
    // rom_array[9597] = 32'h000076f9;
    // rom_array[9598] = 32'h00007701;
    // rom_array[9599] = 32'h00007709;
    // rom_array[9600] = 32'h00007711;
    // rom_array[9601] = 32'h00007719;
    // rom_array[9602] = 32'h00007721;
    // rom_array[9603] = 32'h00007729;
    // rom_array[9604] = 32'h00007731;
    // rom_array[9605] = 32'hFFFFFFF1;
    // rom_array[9606] = 32'hFFFFFFF1;
    // rom_array[9607] = 32'hFFFFFFF1;
    // rom_array[9608] = 32'hFFFFFFF1;
    // rom_array[9609] = 32'h00007739;
    // rom_array[9610] = 32'h00007741;
    // rom_array[9611] = 32'h00007749;
    // rom_array[9612] = 32'h00007751;
    // rom_array[9613] = 32'h00007759;
    // rom_array[9614] = 32'h00007761;
    // rom_array[9615] = 32'h00007769;
    // rom_array[9616] = 32'h00007771;
    // rom_array[9617] = 32'hFFFFFFF0;
    // rom_array[9618] = 32'hFFFFFFF0;
    // rom_array[9619] = 32'hFFFFFFF0;
    // rom_array[9620] = 32'hFFFFFFF0;
    // rom_array[9621] = 32'h00007779;
    // rom_array[9622] = 32'h00007781;
    // rom_array[9623] = 32'hFFFFFFF0;
    // rom_array[9624] = 32'hFFFFFFF0;
    // rom_array[9625] = 32'h00007789;
    // rom_array[9626] = 32'h00007791;
    // rom_array[9627] = 32'h00007799;
    // rom_array[9628] = 32'h000077a1;
    // rom_array[9629] = 32'h000077a9;
    // rom_array[9630] = 32'h000077b1;
    // rom_array[9631] = 32'h000077b9;
    // rom_array[9632] = 32'h000077c1;
    // rom_array[9633] = 32'h000077c9;
    // rom_array[9634] = 32'h000077d1;
    // rom_array[9635] = 32'hFFFFFFF0;
    // rom_array[9636] = 32'hFFFFFFF0;
    // rom_array[9637] = 32'h000077d9;
    // rom_array[9638] = 32'h000077e1;
    // rom_array[9639] = 32'hFFFFFFF0;
    // rom_array[9640] = 32'hFFFFFFF0;
    // rom_array[9641] = 32'h000077e9;
    // rom_array[9642] = 32'h000077f1;
    // rom_array[9643] = 32'h000077f9;
    // rom_array[9644] = 32'h00007801;
    // rom_array[9645] = 32'hFFFFFFF1;
    // rom_array[9646] = 32'hFFFFFFF1;
    // rom_array[9647] = 32'hFFFFFFF1;
    // rom_array[9648] = 32'hFFFFFFF1;
    // rom_array[9649] = 32'h00007809;
    // rom_array[9650] = 32'h00007811;
    // rom_array[9651] = 32'h00007819;
    // rom_array[9652] = 32'h00007821;
    // rom_array[9653] = 32'hFFFFFFF1;
    // rom_array[9654] = 32'hFFFFFFF1;
    // rom_array[9655] = 32'hFFFFFFF1;
    // rom_array[9656] = 32'hFFFFFFF1;
    // rom_array[9657] = 32'h00007829;
    // rom_array[9658] = 32'h00007831;
    // rom_array[9659] = 32'hFFFFFFF1;
    // rom_array[9660] = 32'hFFFFFFF1;
    // rom_array[9661] = 32'h00007839;
    // rom_array[9662] = 32'h00007841;
    // rom_array[9663] = 32'hFFFFFFF1;
    // rom_array[9664] = 32'hFFFFFFF1;
    // rom_array[9665] = 32'h00007849;
    // rom_array[9666] = 32'h00007851;
    // rom_array[9667] = 32'h00007859;
    // rom_array[9668] = 32'h00007861;
    // rom_array[9669] = 32'h00007869;
    // rom_array[9670] = 32'h00007871;
    // rom_array[9671] = 32'hFFFFFFF1;
    // rom_array[9672] = 32'hFFFFFFF1;
    // rom_array[9673] = 32'h00007879;
    // rom_array[9674] = 32'h00007881;
    // rom_array[9675] = 32'h00007889;
    // rom_array[9676] = 32'h00007891;
    // rom_array[9677] = 32'hFFFFFFF1;
    // rom_array[9678] = 32'hFFFFFFF1;
    // rom_array[9679] = 32'h00007899;
    // rom_array[9680] = 32'h000078a1;
    // rom_array[9681] = 32'h000078a9;
    // rom_array[9682] = 32'h000078b1;
    // rom_array[9683] = 32'hFFFFFFF1;
    // rom_array[9684] = 32'hFFFFFFF1;
    // rom_array[9685] = 32'h000078b9;
    // rom_array[9686] = 32'h000078c1;
    // rom_array[9687] = 32'hFFFFFFF1;
    // rom_array[9688] = 32'hFFFFFFF1;
    // rom_array[9689] = 32'hFFFFFFF1;
    // rom_array[9690] = 32'hFFFFFFF1;
    // rom_array[9691] = 32'h000078c9;
    // rom_array[9692] = 32'h000078d1;
    // rom_array[9693] = 32'hFFFFFFF1;
    // rom_array[9694] = 32'hFFFFFFF1;
    // rom_array[9695] = 32'h000078d9;
    // rom_array[9696] = 32'h000078e1;
    // rom_array[9697] = 32'h000078e9;
    // rom_array[9698] = 32'h000078f1;
    // rom_array[9699] = 32'h000078f9;
    // rom_array[9700] = 32'h00007901;
    // rom_array[9701] = 32'hFFFFFFF0;
    // rom_array[9702] = 32'hFFFFFFF0;
    // rom_array[9703] = 32'hFFFFFFF0;
    // rom_array[9704] = 32'hFFFFFFF0;
    // rom_array[9705] = 32'h00007909;
    // rom_array[9706] = 32'h00007911;
    // rom_array[9707] = 32'h00007919;
    // rom_array[9708] = 32'h00007921;
    // rom_array[9709] = 32'hFFFFFFF1;
    // rom_array[9710] = 32'hFFFFFFF1;
    // rom_array[9711] = 32'h00007929;
    // rom_array[9712] = 32'h00007931;
    // rom_array[9713] = 32'h00007939;
    // rom_array[9714] = 32'h00007941;
    // rom_array[9715] = 32'h00007949;
    // rom_array[9716] = 32'h00007951;
    // rom_array[9717] = 32'h00007959;
    // rom_array[9718] = 32'h00007961;
    // rom_array[9719] = 32'h00007969;
    // rom_array[9720] = 32'h00007971;
    // rom_array[9721] = 32'h00007979;
    // rom_array[9722] = 32'h00007981;
    // rom_array[9723] = 32'hFFFFFFF1;
    // rom_array[9724] = 32'hFFFFFFF1;
    // rom_array[9725] = 32'h00007989;
    // rom_array[9726] = 32'h00007991;
    // rom_array[9727] = 32'h00007999;
    // rom_array[9728] = 32'h000079a1;
    // rom_array[9729] = 32'hFFFFFFF1;
    // rom_array[9730] = 32'hFFFFFFF1;
    // rom_array[9731] = 32'hFFFFFFF1;
    // rom_array[9732] = 32'hFFFFFFF1;
    // rom_array[9733] = 32'h000079a9;
    // rom_array[9734] = 32'h000079b1;
    // rom_array[9735] = 32'h000079b9;
    // rom_array[9736] = 32'h000079c1;
    // rom_array[9737] = 32'hFFFFFFF1;
    // rom_array[9738] = 32'hFFFFFFF1;
    // rom_array[9739] = 32'hFFFFFFF1;
    // rom_array[9740] = 32'hFFFFFFF1;
    // rom_array[9741] = 32'h000079c9;
    // rom_array[9742] = 32'h000079d1;
    // rom_array[9743] = 32'h000079d9;
    // rom_array[9744] = 32'h000079e1;
    // rom_array[9745] = 32'hFFFFFFF1;
    // rom_array[9746] = 32'hFFFFFFF1;
    // rom_array[9747] = 32'hFFFFFFF1;
    // rom_array[9748] = 32'hFFFFFFF1;
    // rom_array[9749] = 32'h000079e9;
    // rom_array[9750] = 32'h000079f1;
    // rom_array[9751] = 32'h000079f9;
    // rom_array[9752] = 32'h00007a01;
    // rom_array[9753] = 32'hFFFFFFF1;
    // rom_array[9754] = 32'hFFFFFFF1;
    // rom_array[9755] = 32'h00007a09;
    // rom_array[9756] = 32'h00007a11;
    // rom_array[9757] = 32'h00007a19;
    // rom_array[9758] = 32'h00007a21;
    // rom_array[9759] = 32'h00007a29;
    // rom_array[9760] = 32'h00007a31;
    // rom_array[9761] = 32'hFFFFFFF0;
    // rom_array[9762] = 32'hFFFFFFF0;
    // rom_array[9763] = 32'hFFFFFFF0;
    // rom_array[9764] = 32'hFFFFFFF0;
    // rom_array[9765] = 32'h00007a39;
    // rom_array[9766] = 32'h00007a41;
    // rom_array[9767] = 32'h00007a49;
    // rom_array[9768] = 32'h00007a51;
    // rom_array[9769] = 32'hFFFFFFF0;
    // rom_array[9770] = 32'hFFFFFFF0;
    // rom_array[9771] = 32'hFFFFFFF0;
    // rom_array[9772] = 32'hFFFFFFF0;
    // rom_array[9773] = 32'h00007a59;
    // rom_array[9774] = 32'h00007a61;
    // rom_array[9775] = 32'h00007a69;
    // rom_array[9776] = 32'h00007a71;
    // rom_array[9777] = 32'h00007a79;
    // rom_array[9778] = 32'h00007a81;
    // rom_array[9779] = 32'hFFFFFFF1;
    // rom_array[9780] = 32'hFFFFFFF1;
    // rom_array[9781] = 32'h00007a89;
    // rom_array[9782] = 32'h00007a91;
    // rom_array[9783] = 32'hFFFFFFF1;
    // rom_array[9784] = 32'hFFFFFFF1;
    // rom_array[9785] = 32'h00007a99;
    // rom_array[9786] = 32'h00007aa1;
    // rom_array[9787] = 32'hFFFFFFF1;
    // rom_array[9788] = 32'hFFFFFFF1;
    // rom_array[9789] = 32'h00007aa9;
    // rom_array[9790] = 32'h00007ab1;
    // rom_array[9791] = 32'hFFFFFFF1;
    // rom_array[9792] = 32'hFFFFFFF1;
    // rom_array[9793] = 32'h00007ab9;
    // rom_array[9794] = 32'h00007ac1;
    // rom_array[9795] = 32'hFFFFFFF1;
    // rom_array[9796] = 32'hFFFFFFF1;
    // rom_array[9797] = 32'h00007ac9;
    // rom_array[9798] = 32'h00007ad1;
    // rom_array[9799] = 32'hFFFFFFF1;
    // rom_array[9800] = 32'hFFFFFFF1;
    // rom_array[9801] = 32'hFFFFFFF0;
    // rom_array[9802] = 32'hFFFFFFF0;
    // rom_array[9803] = 32'hFFFFFFF0;
    // rom_array[9804] = 32'hFFFFFFF0;
    // rom_array[9805] = 32'h00007ad9;
    // rom_array[9806] = 32'h00007ae1;
    // rom_array[9807] = 32'hFFFFFFF0;
    // rom_array[9808] = 32'hFFFFFFF0;
    // rom_array[9809] = 32'h00007ae9;
    // rom_array[9810] = 32'h00007af1;
    // rom_array[9811] = 32'hFFFFFFF0;
    // rom_array[9812] = 32'hFFFFFFF0;
    // rom_array[9813] = 32'h00007af9;
    // rom_array[9814] = 32'h00007b01;
    // rom_array[9815] = 32'hFFFFFFF0;
    // rom_array[9816] = 32'hFFFFFFF0;
    // rom_array[9817] = 32'h00007b09;
    // rom_array[9818] = 32'h00007b11;
    // rom_array[9819] = 32'hFFFFFFF0;
    // rom_array[9820] = 32'hFFFFFFF0;
    // rom_array[9821] = 32'h00007b19;
    // rom_array[9822] = 32'h00007b21;
    // rom_array[9823] = 32'hFFFFFFF0;
    // rom_array[9824] = 32'hFFFFFFF0;
    // rom_array[9825] = 32'h00007b29;
    // rom_array[9826] = 32'h00007b31;
    // rom_array[9827] = 32'h00007b39;
    // rom_array[9828] = 32'h00007b41;
    // rom_array[9829] = 32'h00007b49;
    // rom_array[9830] = 32'h00007b51;
    // rom_array[9831] = 32'hFFFFFFF1;
    // rom_array[9832] = 32'hFFFFFFF1;
    // rom_array[9833] = 32'h00007b59;
    // rom_array[9834] = 32'h00007b61;
    // rom_array[9835] = 32'h00007b69;
    // rom_array[9836] = 32'h00007b71;
    // rom_array[9837] = 32'hFFFFFFF1;
    // rom_array[9838] = 32'hFFFFFFF1;
    // rom_array[9839] = 32'hFFFFFFF1;
    // rom_array[9840] = 32'hFFFFFFF1;
    // rom_array[9841] = 32'h00007b79;
    // rom_array[9842] = 32'h00007b81;
    // rom_array[9843] = 32'h00007b89;
    // rom_array[9844] = 32'h00007b91;
    // rom_array[9845] = 32'hFFFFFFF1;
    // rom_array[9846] = 32'hFFFFFFF1;
    // rom_array[9847] = 32'hFFFFFFF1;
    // rom_array[9848] = 32'hFFFFFFF1;
    // rom_array[9849] = 32'h00007b99;
    // rom_array[9850] = 32'h00007ba1;
    // rom_array[9851] = 32'h00007ba9;
    // rom_array[9852] = 32'h00007bb1;
    // rom_array[9853] = 32'hFFFFFFF1;
    // rom_array[9854] = 32'hFFFFFFF1;
    // rom_array[9855] = 32'hFFFFFFF1;
    // rom_array[9856] = 32'hFFFFFFF1;
    // rom_array[9857] = 32'h00007bb9;
    // rom_array[9858] = 32'h00007bc1;
    // rom_array[9859] = 32'hFFFFFFF1;
    // rom_array[9860] = 32'hFFFFFFF1;
    // rom_array[9861] = 32'h00007bc9;
    // rom_array[9862] = 32'h00007bd1;
    // rom_array[9863] = 32'hFFFFFFF1;
    // rom_array[9864] = 32'hFFFFFFF1;
    // rom_array[9865] = 32'h00007bd9;
    // rom_array[9866] = 32'h00007be1;
    // rom_array[9867] = 32'hFFFFFFF1;
    // rom_array[9868] = 32'hFFFFFFF1;
    // rom_array[9869] = 32'h00007be9;
    // rom_array[9870] = 32'h00007bf1;
    // rom_array[9871] = 32'hFFFFFFF1;
    // rom_array[9872] = 32'hFFFFFFF1;
    // rom_array[9873] = 32'h00007bf9;
    // rom_array[9874] = 32'h00007c01;
    // rom_array[9875] = 32'hFFFFFFF1;
    // rom_array[9876] = 32'hFFFFFFF1;
    // rom_array[9877] = 32'h00007c09;
    // rom_array[9878] = 32'h00007c11;
    // rom_array[9879] = 32'hFFFFFFF1;
    // rom_array[9880] = 32'hFFFFFFF1;
    // rom_array[9881] = 32'h00007c19;
    // rom_array[9882] = 32'h00007c21;
    // rom_array[9883] = 32'hFFFFFFF1;
    // rom_array[9884] = 32'hFFFFFFF1;
    // rom_array[9885] = 32'h00007c29;
    // rom_array[9886] = 32'h00007c31;
    // rom_array[9887] = 32'h00007c39;
    // rom_array[9888] = 32'h00007c41;
    // rom_array[9889] = 32'hFFFFFFF1;
    // rom_array[9890] = 32'hFFFFFFF1;
    // rom_array[9891] = 32'hFFFFFFF1;
    // rom_array[9892] = 32'hFFFFFFF1;
    // rom_array[9893] = 32'h00007c49;
    // rom_array[9894] = 32'h00007c51;
    // rom_array[9895] = 32'h00007c59;
    // rom_array[9896] = 32'h00007c61;
    // rom_array[9897] = 32'h00007c69;
    // rom_array[9898] = 32'h00007c71;
    // rom_array[9899] = 32'hFFFFFFF1;
    // rom_array[9900] = 32'hFFFFFFF1;
    // rom_array[9901] = 32'h00007c79;
    // rom_array[9902] = 32'h00007c81;
    // rom_array[9903] = 32'hFFFFFFF1;
    // rom_array[9904] = 32'hFFFFFFF1;
    // rom_array[9905] = 32'h00007c89;
    // rom_array[9906] = 32'h00007c91;
    // rom_array[9907] = 32'h00007c99;
    // rom_array[9908] = 32'h00007ca1;
    // rom_array[9909] = 32'h00007ca9;
    // rom_array[9910] = 32'h00007cb1;
    // rom_array[9911] = 32'hFFFFFFF0;
    // rom_array[9912] = 32'hFFFFFFF0;
    // rom_array[9913] = 32'h00007cb9;
    // rom_array[9914] = 32'h00007cc1;
    // rom_array[9915] = 32'h00007cc9;
    // rom_array[9916] = 32'h00007cd1;
    // rom_array[9917] = 32'hFFFFFFF0;
    // rom_array[9918] = 32'hFFFFFFF0;
    // rom_array[9919] = 32'hFFFFFFF0;
    // rom_array[9920] = 32'hFFFFFFF0;
    // rom_array[9921] = 32'h00007cd9;
    // rom_array[9922] = 32'h00007ce1;
    // rom_array[9923] = 32'h00007ce9;
    // rom_array[9924] = 32'h00007cf1;
    // rom_array[9925] = 32'hFFFFFFF0;
    // rom_array[9926] = 32'hFFFFFFF0;
    // rom_array[9927] = 32'hFFFFFFF0;
    // rom_array[9928] = 32'hFFFFFFF0;
    // rom_array[9929] = 32'h00007cf9;
    // rom_array[9930] = 32'h00007d01;
    // rom_array[9931] = 32'h00007d09;
    // rom_array[9932] = 32'h00007d11;
    // rom_array[9933] = 32'hFFFFFFF0;
    // rom_array[9934] = 32'hFFFFFFF0;
    // rom_array[9935] = 32'hFFFFFFF0;
    // rom_array[9936] = 32'hFFFFFFF0;
    // rom_array[9937] = 32'h00007d19;
    // rom_array[9938] = 32'h00007d21;
    // rom_array[9939] = 32'hFFFFFFF0;
    // rom_array[9940] = 32'hFFFFFFF0;
    // rom_array[9941] = 32'h00007d29;
    // rom_array[9942] = 32'h00007d31;
    // rom_array[9943] = 32'hFFFFFFF0;
    // rom_array[9944] = 32'hFFFFFFF0;
    // rom_array[9945] = 32'h00007d39;
    // rom_array[9946] = 32'h00007d41;
    // rom_array[9947] = 32'hFFFFFFF0;
    // rom_array[9948] = 32'hFFFFFFF0;
    // rom_array[9949] = 32'h00007d49;
    // rom_array[9950] = 32'h00007d51;
    // rom_array[9951] = 32'hFFFFFFF0;
    // rom_array[9952] = 32'hFFFFFFF0;
    // rom_array[9953] = 32'h00007d59;
    // rom_array[9954] = 32'h00007d61;
    // rom_array[9955] = 32'h00007d69;
    // rom_array[9956] = 32'h00007d71;
    // rom_array[9957] = 32'h00007d79;
    // rom_array[9958] = 32'h00007d81;
    // rom_array[9959] = 32'h00007d89;
    // rom_array[9960] = 32'h00007d91;
    // rom_array[9961] = 32'h00007d99;
    // rom_array[9962] = 32'h00007da1;
    // rom_array[9963] = 32'h00007da9;
    // rom_array[9964] = 32'h00007db1;
    // rom_array[9965] = 32'h00007db9;
    // rom_array[9966] = 32'h00007dc1;
    // rom_array[9967] = 32'hFFFFFFF1;
    // rom_array[9968] = 32'hFFFFFFF1;
    // rom_array[9969] = 32'h00007dc9;
    // rom_array[9970] = 32'h00007dd1;
    // rom_array[9971] = 32'hFFFFFFF1;
    // rom_array[9972] = 32'hFFFFFFF1;
    // rom_array[9973] = 32'h00007dd9;
    // rom_array[9974] = 32'h00007de1;
    // rom_array[9975] = 32'h00007de9;
    // rom_array[9976] = 32'h00007df1;
    // rom_array[9977] = 32'h00007df9;
    // rom_array[9978] = 32'h00007e01;
    // rom_array[9979] = 32'hFFFFFFF0;
    // rom_array[9980] = 32'hFFFFFFF0;
    // rom_array[9981] = 32'h00007e09;
    // rom_array[9982] = 32'h00007e11;
    // rom_array[9983] = 32'hFFFFFFF0;
    // rom_array[9984] = 32'hFFFFFFF0;
    // rom_array[9985] = 32'h00007e19;
    // rom_array[9986] = 32'h00007e21;
    // rom_array[9987] = 32'h00007e29;
    // rom_array[9988] = 32'h00007e31;
    // rom_array[9989] = 32'h00007e39;
    // rom_array[9990] = 32'h00007e41;
    // rom_array[9991] = 32'hFFFFFFF1;
    // rom_array[9992] = 32'hFFFFFFF1;
    // rom_array[9993] = 32'h00007e49;
    // rom_array[9994] = 32'h00007e51;
    // rom_array[9995] = 32'hFFFFFFF0;
    // rom_array[9996] = 32'hFFFFFFF0;
    // rom_array[9997] = 32'hFFFFFFF0;
    // rom_array[9998] = 32'hFFFFFFF0;
    // rom_array[9999] = 32'hFFFFFFF0;
    // rom_array[10000] = 32'hFFFFFFF0;
    // rom_array[10001] = 32'h00007e59;
    // rom_array[10002] = 32'h00007e61;
    // rom_array[10003] = 32'hFFFFFFF1;
    // rom_array[10004] = 32'hFFFFFFF1;
    // rom_array[10005] = 32'h00007e69;
    // rom_array[10006] = 32'h00007e71;
    // rom_array[10007] = 32'hFFFFFFF1;
    // rom_array[10008] = 32'hFFFFFFF1;
    // rom_array[10009] = 32'h00007e79;
    // rom_array[10010] = 32'h00007e81;
    // rom_array[10011] = 32'h00007e89;
    // rom_array[10012] = 32'h00007e91;
    // rom_array[10013] = 32'hFFFFFFF1;
    // rom_array[10014] = 32'hFFFFFFF1;
    // rom_array[10015] = 32'hFFFFFFF1;
    // rom_array[10016] = 32'hFFFFFFF1;
    // rom_array[10017] = 32'h00007e99;
    // rom_array[10018] = 32'h00007ea1;
    // rom_array[10019] = 32'h00007ea9;
    // rom_array[10020] = 32'h00007eb1;
    // rom_array[10021] = 32'hFFFFFFF1;
    // rom_array[10022] = 32'hFFFFFFF1;
    // rom_array[10023] = 32'hFFFFFFF1;
    // rom_array[10024] = 32'hFFFFFFF1;
    // rom_array[10025] = 32'h00007eb9;
    // rom_array[10026] = 32'h00007ec1;
    // rom_array[10027] = 32'h00007ec9;
    // rom_array[10028] = 32'h00007ed1;
    // rom_array[10029] = 32'hFFFFFFF1;
    // rom_array[10030] = 32'hFFFFFFF1;
    // rom_array[10031] = 32'hFFFFFFF1;
    // rom_array[10032] = 32'hFFFFFFF1;
    // rom_array[10033] = 32'h00007ed9;
    // rom_array[10034] = 32'h00007ee1;
    // rom_array[10035] = 32'h00007ee9;
    // rom_array[10036] = 32'h00007ef1;
    // rom_array[10037] = 32'hFFFFFFF1;
    // rom_array[10038] = 32'hFFFFFFF1;
    // rom_array[10039] = 32'hFFFFFFF1;
    // rom_array[10040] = 32'hFFFFFFF1;
    // rom_array[10041] = 32'hFFFFFFF0;
    // rom_array[10042] = 32'hFFFFFFF0;
    // rom_array[10043] = 32'hFFFFFFF0;
    // rom_array[10044] = 32'hFFFFFFF0;
    // rom_array[10045] = 32'h00007ef9;
    // rom_array[10046] = 32'h00007f01;
    // rom_array[10047] = 32'h00007f09;
    // rom_array[10048] = 32'h00007f11;
    // rom_array[10049] = 32'hFFFFFFF0;
    // rom_array[10050] = 32'hFFFFFFF0;
    // rom_array[10051] = 32'hFFFFFFF0;
    // rom_array[10052] = 32'hFFFFFFF0;
    // rom_array[10053] = 32'h00007f19;
    // rom_array[10054] = 32'h00007f21;
    // rom_array[10055] = 32'h00007f29;
    // rom_array[10056] = 32'h00007f31;
    // rom_array[10057] = 32'h00007f39;
    // rom_array[10058] = 32'h00007f41;
    // rom_array[10059] = 32'hFFFFFFF1;
    // rom_array[10060] = 32'hFFFFFFF1;
    // rom_array[10061] = 32'h00007f49;
    // rom_array[10062] = 32'h00007f51;
    // rom_array[10063] = 32'hFFFFFFF1;
    // rom_array[10064] = 32'hFFFFFFF1;
    // rom_array[10065] = 32'hFFFFFFF0;
    // rom_array[10066] = 32'hFFFFFFF0;
    // rom_array[10067] = 32'hFFFFFFF0;
    // rom_array[10068] = 32'hFFFFFFF0;
    // rom_array[10069] = 32'h00007f59;
    // rom_array[10070] = 32'h00007f61;
    // rom_array[10071] = 32'hFFFFFFF0;
    // rom_array[10072] = 32'hFFFFFFF0;
    // rom_array[10073] = 32'h00007f69;
    // rom_array[10074] = 32'h00007f71;
    // rom_array[10075] = 32'hFFFFFFF0;
    // rom_array[10076] = 32'hFFFFFFF0;
    // rom_array[10077] = 32'h00007f79;
    // rom_array[10078] = 32'h00007f81;
    // rom_array[10079] = 32'hFFFFFFF0;
    // rom_array[10080] = 32'hFFFFFFF0;
    // rom_array[10081] = 32'h00007f89;
    // rom_array[10082] = 32'h00007f91;
    // rom_array[10083] = 32'h00007f99;
    // rom_array[10084] = 32'h00007fa1;
    // rom_array[10085] = 32'h00007fa9;
    // rom_array[10086] = 32'h00007fb1;
    // rom_array[10087] = 32'hFFFFFFF1;
    // rom_array[10088] = 32'hFFFFFFF1;
    // rom_array[10089] = 32'h00007fb9;
    // rom_array[10090] = 32'h00007fc1;
    // rom_array[10091] = 32'h00007fc9;
    // rom_array[10092] = 32'h00007fd1;
    // rom_array[10093] = 32'hFFFFFFF1;
    // rom_array[10094] = 32'hFFFFFFF1;
    // rom_array[10095] = 32'hFFFFFFF1;
    // rom_array[10096] = 32'hFFFFFFF1;
    // rom_array[10097] = 32'h00007fd9;
    // rom_array[10098] = 32'h00007fe1;
    // rom_array[10099] = 32'hFFFFFFF1;
    // rom_array[10100] = 32'hFFFFFFF1;
    // rom_array[10101] = 32'h00007fe9;
    // rom_array[10102] = 32'h00007ff1;
    // rom_array[10103] = 32'hFFFFFFF1;
    // rom_array[10104] = 32'hFFFFFFF1;
    // rom_array[10105] = 32'h00007ff9;
    // rom_array[10106] = 32'h00008001;
    // rom_array[10107] = 32'h00008009;
    // rom_array[10108] = 32'h00008011;
    // rom_array[10109] = 32'h00008019;
    // rom_array[10110] = 32'h00008021;
    // rom_array[10111] = 32'hFFFFFFF1;
    // rom_array[10112] = 32'hFFFFFFF1;
    // rom_array[10113] = 32'h00008029;
    // rom_array[10114] = 32'h00008031;
    // rom_array[10115] = 32'h00008039;
    // rom_array[10116] = 32'h00008041;
    // rom_array[10117] = 32'hFFFFFFF0;
    // rom_array[10118] = 32'hFFFFFFF0;
    // rom_array[10119] = 32'hFFFFFFF0;
    // rom_array[10120] = 32'hFFFFFFF0;
    // rom_array[10121] = 32'h00008049;
    // rom_array[10122] = 32'h00008051;
    // rom_array[10123] = 32'hFFFFFFF1;
    // rom_array[10124] = 32'hFFFFFFF1;
    // rom_array[10125] = 32'h00008059;
    // rom_array[10126] = 32'h00008061;
    // rom_array[10127] = 32'hFFFFFFF1;
    // rom_array[10128] = 32'hFFFFFFF1;
    // rom_array[10129] = 32'h00008069;
    // rom_array[10130] = 32'h00008071;
    // rom_array[10131] = 32'h00008079;
    // rom_array[10132] = 32'h00008081;
    // rom_array[10133] = 32'h00008089;
    // rom_array[10134] = 32'h00008091;
    // rom_array[10135] = 32'hFFFFFFF1;
    // rom_array[10136] = 32'hFFFFFFF1;
    // rom_array[10137] = 32'h00008099;
    // rom_array[10138] = 32'h000080a1;
    // rom_array[10139] = 32'h000080a9;
    // rom_array[10140] = 32'h000080b1;
    // rom_array[10141] = 32'hFFFFFFF1;
    // rom_array[10142] = 32'hFFFFFFF1;
    // rom_array[10143] = 32'hFFFFFFF1;
    // rom_array[10144] = 32'hFFFFFFF1;
    // rom_array[10145] = 32'h000080b9;
    // rom_array[10146] = 32'h000080c1;
    // rom_array[10147] = 32'hFFFFFFF1;
    // rom_array[10148] = 32'hFFFFFFF1;
    // rom_array[10149] = 32'h000080c9;
    // rom_array[10150] = 32'h000080d1;
    // rom_array[10151] = 32'hFFFFFFF1;
    // rom_array[10152] = 32'hFFFFFFF1;
    // rom_array[10153] = 32'h000080d9;
    // rom_array[10154] = 32'h000080e1;
    // rom_array[10155] = 32'h000080e9;
    // rom_array[10156] = 32'h000080f1;
    // rom_array[10157] = 32'h000080f9;
    // rom_array[10158] = 32'h00008101;
    // rom_array[10159] = 32'hFFFFFFF1;
    // rom_array[10160] = 32'hFFFFFFF1;
    // rom_array[10161] = 32'h00008109;
    // rom_array[10162] = 32'h00008111;
    // rom_array[10163] = 32'h00008119;
    // rom_array[10164] = 32'h00008121;
    // rom_array[10165] = 32'hFFFFFFF1;
    // rom_array[10166] = 32'hFFFFFFF1;
    // rom_array[10167] = 32'hFFFFFFF1;
    // rom_array[10168] = 32'hFFFFFFF1;
    // rom_array[10169] = 32'h00008129;
    // rom_array[10170] = 32'h00008131;
    // rom_array[10171] = 32'hFFFFFFF0;
    // rom_array[10172] = 32'hFFFFFFF0;
    // rom_array[10173] = 32'h00008139;
    // rom_array[10174] = 32'h00008141;
    // rom_array[10175] = 32'hFFFFFFF0;
    // rom_array[10176] = 32'hFFFFFFF0;
    // rom_array[10177] = 32'h00008149;
    // rom_array[10178] = 32'h00008151;
    // rom_array[10179] = 32'h00008159;
    // rom_array[10180] = 32'h00008161;
    // rom_array[10181] = 32'h00008169;
    // rom_array[10182] = 32'h00008171;
    // rom_array[10183] = 32'hFFFFFFF1;
    // rom_array[10184] = 32'hFFFFFFF1;
    // rom_array[10185] = 32'h00008179;
    // rom_array[10186] = 32'h00008181;
    // rom_array[10187] = 32'h00008189;
    // rom_array[10188] = 32'h00008191;
    // rom_array[10189] = 32'hFFFFFFF0;
    // rom_array[10190] = 32'hFFFFFFF0;
    // rom_array[10191] = 32'hFFFFFFF0;
    // rom_array[10192] = 32'hFFFFFFF0;
    // rom_array[10193] = 32'h00008199;
    // rom_array[10194] = 32'h000081a1;
    // rom_array[10195] = 32'hFFFFFFF1;
    // rom_array[10196] = 32'hFFFFFFF1;
    // rom_array[10197] = 32'h000081a9;
    // rom_array[10198] = 32'h000081b1;
    // rom_array[10199] = 32'h000081b9;
    // rom_array[10200] = 32'h000081c1;
    // rom_array[10201] = 32'hFFFFFFF1;
    // rom_array[10202] = 32'hFFFFFFF1;
    // rom_array[10203] = 32'hFFFFFFF1;
    // rom_array[10204] = 32'hFFFFFFF1;
    // rom_array[10205] = 32'h000081c9;
    // rom_array[10206] = 32'h000081d1;
    // rom_array[10207] = 32'h000081d9;
    // rom_array[10208] = 32'h000081e1;
    // rom_array[10209] = 32'h000081e9;
    // rom_array[10210] = 32'h000081f1;
    // rom_array[10211] = 32'h000081f9;
    // rom_array[10212] = 32'h00008201;
    // rom_array[10213] = 32'h00008209;
    // rom_array[10214] = 32'h00008211;
    // rom_array[10215] = 32'hFFFFFFF0;
    // rom_array[10216] = 32'hFFFFFFF0;
    // rom_array[10217] = 32'h00008219;
    // rom_array[10218] = 32'h00008221;
    // rom_array[10219] = 32'h00008229;
    // rom_array[10220] = 32'h00008231;
    // rom_array[10221] = 32'hFFFFFFF0;
    // rom_array[10222] = 32'hFFFFFFF0;
    // rom_array[10223] = 32'hFFFFFFF0;
    // rom_array[10224] = 32'hFFFFFFF0;
    // rom_array[10225] = 32'h00008239;
    // rom_array[10226] = 32'h00008241;
    // rom_array[10227] = 32'hFFFFFFF0;
    // rom_array[10228] = 32'hFFFFFFF0;
    // rom_array[10229] = 32'h00008249;
    // rom_array[10230] = 32'h00008251;
    // rom_array[10231] = 32'hFFFFFFF0;
    // rom_array[10232] = 32'hFFFFFFF0;
    // rom_array[10233] = 32'h00008259;
    // rom_array[10234] = 32'h00008261;
    // rom_array[10235] = 32'h00008269;
    // rom_array[10236] = 32'h00008271;
    // rom_array[10237] = 32'h00008279;
    // rom_array[10238] = 32'h00008281;
    // rom_array[10239] = 32'h00008289;
    // rom_array[10240] = 32'h00008291;
    // rom_array[10241] = 32'h00008299;
    // rom_array[10242] = 32'h000082a1;
    // rom_array[10243] = 32'hFFFFFFF0;
    // rom_array[10244] = 32'hFFFFFFF0;
    // rom_array[10245] = 32'h000082a9;
    // rom_array[10246] = 32'h000082b1;
    // rom_array[10247] = 32'hFFFFFFF0;
    // rom_array[10248] = 32'hFFFFFFF0;
    // rom_array[10249] = 32'h000082b9;
    // rom_array[10250] = 32'h000082c1;
    // rom_array[10251] = 32'hFFFFFFF1;
    // rom_array[10252] = 32'hFFFFFFF1;
    // rom_array[10253] = 32'h000082c9;
    // rom_array[10254] = 32'h000082d1;
    // rom_array[10255] = 32'h000082d9;
    // rom_array[10256] = 32'h000082e1;
    // rom_array[10257] = 32'h000082e9;
    // rom_array[10258] = 32'h000082f1;
    // rom_array[10259] = 32'hFFFFFFF0;
    // rom_array[10260] = 32'hFFFFFFF0;
    // rom_array[10261] = 32'h000082f9;
    // rom_array[10262] = 32'h00008301;
    // rom_array[10263] = 32'hFFFFFFF0;
    // rom_array[10264] = 32'hFFFFFFF0;
    // rom_array[10265] = 32'h00008309;
    // rom_array[10266] = 32'h00008311;
    // rom_array[10267] = 32'h00008319;
    // rom_array[10268] = 32'h00008321;
    // rom_array[10269] = 32'hFFFFFFF0;
    // rom_array[10270] = 32'hFFFFFFF0;
    // rom_array[10271] = 32'hFFFFFFF0;
    // rom_array[10272] = 32'hFFFFFFF0;
    // rom_array[10273] = 32'h00008329;
    // rom_array[10274] = 32'h00008331;
    // rom_array[10275] = 32'h00008339;
    // rom_array[10276] = 32'h00008341;
    // rom_array[10277] = 32'hFFFFFFF0;
    // rom_array[10278] = 32'hFFFFFFF0;
    // rom_array[10279] = 32'hFFFFFFF0;
    // rom_array[10280] = 32'hFFFFFFF0;
    // rom_array[10281] = 32'h00008349;
    // rom_array[10282] = 32'h00008351;
    // rom_array[10283] = 32'h00008359;
    // rom_array[10284] = 32'h00008361;
    // rom_array[10285] = 32'hFFFFFFF0;
    // rom_array[10286] = 32'hFFFFFFF0;
    // rom_array[10287] = 32'hFFFFFFF0;
    // rom_array[10288] = 32'hFFFFFFF0;
    // rom_array[10289] = 32'h00008369;
    // rom_array[10290] = 32'h00008371;
    // rom_array[10291] = 32'h00008379;
    // rom_array[10292] = 32'h00008381;
    // rom_array[10293] = 32'hFFFFFFF0;
    // rom_array[10294] = 32'hFFFFFFF0;
    // rom_array[10295] = 32'hFFFFFFF0;
    // rom_array[10296] = 32'hFFFFFFF0;
    // rom_array[10297] = 32'h00008389;
    // rom_array[10298] = 32'h00008391;
    // rom_array[10299] = 32'h00008399;
    // rom_array[10300] = 32'h000083a1;
    // rom_array[10301] = 32'hFFFFFFF0;
    // rom_array[10302] = 32'hFFFFFFF0;
    // rom_array[10303] = 32'hFFFFFFF0;
    // rom_array[10304] = 32'hFFFFFFF0;
    // rom_array[10305] = 32'h000083a9;
    // rom_array[10306] = 32'h000083b1;
    // rom_array[10307] = 32'h000083b9;
    // rom_array[10308] = 32'h000083c1;
    // rom_array[10309] = 32'hFFFFFFF0;
    // rom_array[10310] = 32'hFFFFFFF0;
    // rom_array[10311] = 32'hFFFFFFF0;
    // rom_array[10312] = 32'hFFFFFFF0;
    // rom_array[10313] = 32'h000083c9;
    // rom_array[10314] = 32'h000083d1;
    // rom_array[10315] = 32'h000083d9;
    // rom_array[10316] = 32'h000083e1;
    // rom_array[10317] = 32'h000083e9;
    // rom_array[10318] = 32'h000083f1;
    // rom_array[10319] = 32'hFFFFFFF1;
    // rom_array[10320] = 32'hFFFFFFF1;
    // rom_array[10321] = 32'h000083f9;
    // rom_array[10322] = 32'h00008401;
    // rom_array[10323] = 32'h00008409;
    // rom_array[10324] = 32'h00008411;
    // rom_array[10325] = 32'hFFFFFFF1;
    // rom_array[10326] = 32'hFFFFFFF1;
    // rom_array[10327] = 32'hFFFFFFF1;
    // rom_array[10328] = 32'hFFFFFFF1;
    // rom_array[10329] = 32'h00008419;
    // rom_array[10330] = 32'h00008421;
    // rom_array[10331] = 32'hFFFFFFF1;
    // rom_array[10332] = 32'hFFFFFFF1;
    // rom_array[10333] = 32'h00008429;
    // rom_array[10334] = 32'h00008431;
    // rom_array[10335] = 32'hFFFFFFF1;
    // rom_array[10336] = 32'hFFFFFFF1;
    // rom_array[10337] = 32'h00008439;
    // rom_array[10338] = 32'h00008441;
    // rom_array[10339] = 32'h00008449;
    // rom_array[10340] = 32'h00008451;
    // rom_array[10341] = 32'hFFFFFFF1;
    // rom_array[10342] = 32'hFFFFFFF1;
    // rom_array[10343] = 32'hFFFFFFF1;
    // rom_array[10344] = 32'hFFFFFFF1;
    // rom_array[10345] = 32'h00008459;
    // rom_array[10346] = 32'h00008461;
    // rom_array[10347] = 32'h00008469;
    // rom_array[10348] = 32'h00008471;
    // rom_array[10349] = 32'hFFFFFFF1;
    // rom_array[10350] = 32'hFFFFFFF1;
    // rom_array[10351] = 32'hFFFFFFF1;
    // rom_array[10352] = 32'hFFFFFFF1;
    // rom_array[10353] = 32'h00008479;
    // rom_array[10354] = 32'h00008481;
    // rom_array[10355] = 32'h00008489;
    // rom_array[10356] = 32'h00008491;
    // rom_array[10357] = 32'hFFFFFFF1;
    // rom_array[10358] = 32'hFFFFFFF1;
    // rom_array[10359] = 32'hFFFFFFF1;
    // rom_array[10360] = 32'hFFFFFFF1;
    // rom_array[10361] = 32'h00008499;
    // rom_array[10362] = 32'h000084a1;
    // rom_array[10363] = 32'h000084a9;
    // rom_array[10364] = 32'h000084b1;
    // rom_array[10365] = 32'hFFFFFFF1;
    // rom_array[10366] = 32'hFFFFFFF1;
    // rom_array[10367] = 32'hFFFFFFF1;
    // rom_array[10368] = 32'hFFFFFFF1;
    // rom_array[10369] = 32'h000084b9;
    // rom_array[10370] = 32'h000084c1;
    // rom_array[10371] = 32'h000084c9;
    // rom_array[10372] = 32'h000084d1;
    // rom_array[10373] = 32'h000084d9;
    // rom_array[10374] = 32'h000084e1;
    // rom_array[10375] = 32'hFFFFFFF1;
    // rom_array[10376] = 32'hFFFFFFF1;
    // rom_array[10377] = 32'h000084e9;
    // rom_array[10378] = 32'h000084f1;
    // rom_array[10379] = 32'h000084f9;
    // rom_array[10380] = 32'h00008501;
    // rom_array[10381] = 32'hFFFFFFF1;
    // rom_array[10382] = 32'hFFFFFFF1;
    // rom_array[10383] = 32'hFFFFFFF1;
    // rom_array[10384] = 32'hFFFFFFF1;
    // rom_array[10385] = 32'h00008509;
    // rom_array[10386] = 32'h00008511;
    // rom_array[10387] = 32'hFFFFFFF1;
    // rom_array[10388] = 32'hFFFFFFF1;
    // rom_array[10389] = 32'h00008519;
    // rom_array[10390] = 32'h00008521;
    // rom_array[10391] = 32'hFFFFFFF1;
    // rom_array[10392] = 32'hFFFFFFF1;
    // rom_array[10393] = 32'h00008529;
    // rom_array[10394] = 32'h00008531;
    // rom_array[10395] = 32'hFFFFFFF1;
    // rom_array[10396] = 32'hFFFFFFF1;
    // rom_array[10397] = 32'h00008539;
    // rom_array[10398] = 32'h00008541;
    // rom_array[10399] = 32'hFFFFFFF1;
    // rom_array[10400] = 32'hFFFFFFF1;
    // rom_array[10401] = 32'h00008549;
    // rom_array[10402] = 32'h00008551;
    // rom_array[10403] = 32'hFFFFFFF1;
    // rom_array[10404] = 32'hFFFFFFF1;
    // rom_array[10405] = 32'h00008559;
    // rom_array[10406] = 32'h00008561;
    // rom_array[10407] = 32'hFFFFFFF1;
    // rom_array[10408] = 32'hFFFFFFF1;
    // rom_array[10409] = 32'h00008569;
    // rom_array[10410] = 32'h00008571;
    // rom_array[10411] = 32'h00008579;
    // rom_array[10412] = 32'h00008581;
    // rom_array[10413] = 32'h00008589;
    // rom_array[10414] = 32'h00008591;
    // rom_array[10415] = 32'hFFFFFFF0;
    // rom_array[10416] = 32'hFFFFFFF0;
    // rom_array[10417] = 32'h00008599;
    // rom_array[10418] = 32'h000085a1;
    // rom_array[10419] = 32'h000085a9;
    // rom_array[10420] = 32'h000085b1;
    // rom_array[10421] = 32'hFFFFFFF0;
    // rom_array[10422] = 32'hFFFFFFF0;
    // rom_array[10423] = 32'hFFFFFFF0;
    // rom_array[10424] = 32'hFFFFFFF0;
    // rom_array[10425] = 32'h000085b9;
    // rom_array[10426] = 32'h000085c1;
    // rom_array[10427] = 32'hFFFFFFF0;
    // rom_array[10428] = 32'hFFFFFFF0;
    // rom_array[10429] = 32'h000085c9;
    // rom_array[10430] = 32'h000085d1;
    // rom_array[10431] = 32'hFFFFFFF0;
    // rom_array[10432] = 32'hFFFFFFF0;
    // rom_array[10433] = 32'h000085d9;
    // rom_array[10434] = 32'h000085e1;
    // rom_array[10435] = 32'h000085e9;
    // rom_array[10436] = 32'h000085f1;
    // rom_array[10437] = 32'hFFFFFFF0;
    // rom_array[10438] = 32'hFFFFFFF0;
    // rom_array[10439] = 32'hFFFFFFF0;
    // rom_array[10440] = 32'hFFFFFFF0;
    // rom_array[10441] = 32'h000085f9;
    // rom_array[10442] = 32'h00008601;
    // rom_array[10443] = 32'h00008609;
    // rom_array[10444] = 32'h00008611;
    // rom_array[10445] = 32'hFFFFFFF0;
    // rom_array[10446] = 32'hFFFFFFF0;
    // rom_array[10447] = 32'hFFFFFFF0;
    // rom_array[10448] = 32'hFFFFFFF0;
    // rom_array[10449] = 32'h00008619;
    // rom_array[10450] = 32'h00008621;
    // rom_array[10451] = 32'hFFFFFFF0;
    // rom_array[10452] = 32'hFFFFFFF0;
    // rom_array[10453] = 32'h00008629;
    // rom_array[10454] = 32'h00008631;
    // rom_array[10455] = 32'hFFFFFFF0;
    // rom_array[10456] = 32'hFFFFFFF0;
    // rom_array[10457] = 32'h00008639;
    // rom_array[10458] = 32'h00008641;
    // rom_array[10459] = 32'hFFFFFFF0;
    // rom_array[10460] = 32'hFFFFFFF0;
    // rom_array[10461] = 32'h00008649;
    // rom_array[10462] = 32'h00008651;
    // rom_array[10463] = 32'hFFFFFFF0;
    // rom_array[10464] = 32'hFFFFFFF0;
    // rom_array[10465] = 32'h00008659;
    // rom_array[10466] = 32'h00008661;
    // rom_array[10467] = 32'hFFFFFFF1;
    // rom_array[10468] = 32'hFFFFFFF1;
    // rom_array[10469] = 32'h00008669;
    // rom_array[10470] = 32'h00008671;
    // rom_array[10471] = 32'hFFFFFFF1;
    // rom_array[10472] = 32'hFFFFFFF1;
    // rom_array[10473] = 32'h00008679;
    // rom_array[10474] = 32'h00008681;
    // rom_array[10475] = 32'h00008689;
    // rom_array[10476] = 32'h00008691;
    // rom_array[10477] = 32'hFFFFFFF0;
    // rom_array[10478] = 32'hFFFFFFF0;
    // rom_array[10479] = 32'hFFFFFFF0;
    // rom_array[10480] = 32'hFFFFFFF0;
    // rom_array[10481] = 32'h00008699;
    // rom_array[10482] = 32'h000086a1;
    // rom_array[10483] = 32'h000086a9;
    // rom_array[10484] = 32'h000086b1;
    // rom_array[10485] = 32'hFFFFFFF0;
    // rom_array[10486] = 32'hFFFFFFF0;
    // rom_array[10487] = 32'hFFFFFFF0;
    // rom_array[10488] = 32'hFFFFFFF0;
    // rom_array[10489] = 32'h000086b9;
    // rom_array[10490] = 32'h000086c1;
    // rom_array[10491] = 32'hFFFFFFF0;
    // rom_array[10492] = 32'hFFFFFFF0;
    // rom_array[10493] = 32'h000086c9;
    // rom_array[10494] = 32'h000086d1;
    // rom_array[10495] = 32'hFFFFFFF0;
    // rom_array[10496] = 32'hFFFFFFF0;
    // rom_array[10497] = 32'h000086d9;
    // rom_array[10498] = 32'h000086e1;
    // rom_array[10499] = 32'hFFFFFFF0;
    // rom_array[10500] = 32'hFFFFFFF0;
    // rom_array[10501] = 32'hFFFFFFF0;
    // rom_array[10502] = 32'hFFFFFFF0;
    // rom_array[10503] = 32'hFFFFFFF0;
    // rom_array[10504] = 32'hFFFFFFF0;
    // rom_array[10505] = 32'h000086e9;
    // rom_array[10506] = 32'h000086f1;
    // rom_array[10507] = 32'h000086f9;
    // rom_array[10508] = 32'h00008701;
    // rom_array[10509] = 32'hFFFFFFF0;
    // rom_array[10510] = 32'hFFFFFFF0;
    // rom_array[10511] = 32'hFFFFFFF0;
    // rom_array[10512] = 32'hFFFFFFF0;
    // rom_array[10513] = 32'h00008709;
    // rom_array[10514] = 32'h00008711;
    // rom_array[10515] = 32'h00008719;
    // rom_array[10516] = 32'h00008721;
    // rom_array[10517] = 32'hFFFFFFF0;
    // rom_array[10518] = 32'hFFFFFFF0;
    // rom_array[10519] = 32'hFFFFFFF0;
    // rom_array[10520] = 32'hFFFFFFF0;
    // rom_array[10521] = 32'h00008729;
    // rom_array[10522] = 32'h00008731;
    // rom_array[10523] = 32'hFFFFFFF0;
    // rom_array[10524] = 32'hFFFFFFF0;
    // rom_array[10525] = 32'hFFFFFFF0;
    // rom_array[10526] = 32'hFFFFFFF0;
    // rom_array[10527] = 32'hFFFFFFF0;
    // rom_array[10528] = 32'hFFFFFFF0;
    // rom_array[10529] = 32'hFFFFFFF0;
    // rom_array[10530] = 32'hFFFFFFF0;
    // rom_array[10531] = 32'h00008739;
    // rom_array[10532] = 32'h00008741;
    // rom_array[10533] = 32'hFFFFFFF0;
    // rom_array[10534] = 32'hFFFFFFF0;
    // rom_array[10535] = 32'hFFFFFFF0;
    // rom_array[10536] = 32'hFFFFFFF0;
    // rom_array[10537] = 32'h00008749;
    // rom_array[10538] = 32'h00008751;
    // rom_array[10539] = 32'h00008759;
    // rom_array[10540] = 32'h00008761;
    // rom_array[10541] = 32'hFFFFFFF0;
    // rom_array[10542] = 32'hFFFFFFF0;
    // rom_array[10543] = 32'hFFFFFFF0;
    // rom_array[10544] = 32'hFFFFFFF0;
    // rom_array[10545] = 32'h00008769;
    // rom_array[10546] = 32'h00008771;
    // rom_array[10547] = 32'h00008779;
    // rom_array[10548] = 32'h00008781;
    // rom_array[10549] = 32'h00008789;
    // rom_array[10550] = 32'h00008791;
    // rom_array[10551] = 32'hFFFFFFF1;
    // rom_array[10552] = 32'hFFFFFFF1;
    // rom_array[10553] = 32'h00008799;
    // rom_array[10554] = 32'h000087a1;
    // rom_array[10555] = 32'h000087a9;
    // rom_array[10556] = 32'h000087b1;
    // rom_array[10557] = 32'hFFFFFFF1;
    // rom_array[10558] = 32'hFFFFFFF1;
    // rom_array[10559] = 32'hFFFFFFF1;
    // rom_array[10560] = 32'hFFFFFFF1;
    // rom_array[10561] = 32'h000087b9;
    // rom_array[10562] = 32'h000087c1;
    // rom_array[10563] = 32'hFFFFFFF1;
    // rom_array[10564] = 32'hFFFFFFF1;
    // rom_array[10565] = 32'h000087c9;
    // rom_array[10566] = 32'h000087d1;
    // rom_array[10567] = 32'hFFFFFFF1;
    // rom_array[10568] = 32'hFFFFFFF1;
    // rom_array[10569] = 32'h000087d9;
    // rom_array[10570] = 32'h000087e1;
    // rom_array[10571] = 32'h000087e9;
    // rom_array[10572] = 32'h000087f1;
    // rom_array[10573] = 32'hFFFFFFF0;
    // rom_array[10574] = 32'hFFFFFFF0;
    // rom_array[10575] = 32'hFFFFFFF0;
    // rom_array[10576] = 32'hFFFFFFF0;
    // rom_array[10577] = 32'h000087f9;
    // rom_array[10578] = 32'h00008801;
    // rom_array[10579] = 32'h00008809;
    // rom_array[10580] = 32'h00008811;
    // rom_array[10581] = 32'hFFFFFFF0;
    // rom_array[10582] = 32'hFFFFFFF0;
    // rom_array[10583] = 32'hFFFFFFF0;
    // rom_array[10584] = 32'hFFFFFFF0;
    // rom_array[10585] = 32'h00008819;
    // rom_array[10586] = 32'h00008821;
    // rom_array[10587] = 32'h00008829;
    // rom_array[10588] = 32'h00008831;
    // rom_array[10589] = 32'hFFFFFFF1;
    // rom_array[10590] = 32'hFFFFFFF1;
    // rom_array[10591] = 32'hFFFFFFF1;
    // rom_array[10592] = 32'hFFFFFFF1;
    // rom_array[10593] = 32'h00008839;
    // rom_array[10594] = 32'h00008841;
    // rom_array[10595] = 32'h00008849;
    // rom_array[10596] = 32'h00008851;
    // rom_array[10597] = 32'hFFFFFFF1;
    // rom_array[10598] = 32'hFFFFFFF1;
    // rom_array[10599] = 32'hFFFFFFF1;
    // rom_array[10600] = 32'hFFFFFFF1;
    // rom_array[10601] = 32'h00008859;
    // rom_array[10602] = 32'h00008861;
    // rom_array[10603] = 32'h00008869;
    // rom_array[10604] = 32'h00008871;
    // rom_array[10605] = 32'hFFFFFFF1;
    // rom_array[10606] = 32'hFFFFFFF1;
    // rom_array[10607] = 32'hFFFFFFF1;
    // rom_array[10608] = 32'hFFFFFFF1;
    // rom_array[10609] = 32'h00008879;
    // rom_array[10610] = 32'h00008881;
    // rom_array[10611] = 32'h00008889;
    // rom_array[10612] = 32'h00008891;
    // rom_array[10613] = 32'hFFFFFFF1;
    // rom_array[10614] = 32'hFFFFFFF1;
    // rom_array[10615] = 32'hFFFFFFF1;
    // rom_array[10616] = 32'hFFFFFFF1;
    // rom_array[10617] = 32'h00008899;
    // rom_array[10618] = 32'h000088a1;
    // rom_array[10619] = 32'h000088a9;
    // rom_array[10620] = 32'h000088b1;
    // rom_array[10621] = 32'hFFFFFFF0;
    // rom_array[10622] = 32'hFFFFFFF0;
    // rom_array[10623] = 32'hFFFFFFF0;
    // rom_array[10624] = 32'hFFFFFFF0;
    // rom_array[10625] = 32'h000088b9;
    // rom_array[10626] = 32'h000088c1;
    // rom_array[10627] = 32'h000088c9;
    // rom_array[10628] = 32'h000088d1;
    // rom_array[10629] = 32'hFFFFFFF0;
    // rom_array[10630] = 32'hFFFFFFF0;
    // rom_array[10631] = 32'hFFFFFFF0;
    // rom_array[10632] = 32'hFFFFFFF0;
    // rom_array[10633] = 32'h000088d9;
    // rom_array[10634] = 32'h000088e1;
    // rom_array[10635] = 32'h000088e9;
    // rom_array[10636] = 32'h000088f1;
    // rom_array[10637] = 32'h000088f9;
    // rom_array[10638] = 32'h00008901;
    // rom_array[10639] = 32'hFFFFFFF1;
    // rom_array[10640] = 32'hFFFFFFF1;
    // rom_array[10641] = 32'h00008909;
    // rom_array[10642] = 32'h00008911;
    // rom_array[10643] = 32'h00008919;
    // rom_array[10644] = 32'h00008921;
    // rom_array[10645] = 32'hFFFFFFF1;
    // rom_array[10646] = 32'hFFFFFFF1;
    // rom_array[10647] = 32'hFFFFFFF1;
    // rom_array[10648] = 32'hFFFFFFF1;
    // rom_array[10649] = 32'h00008929;
    // rom_array[10650] = 32'h00008931;
    // rom_array[10651] = 32'h00008939;
    // rom_array[10652] = 32'h00008941;
    // rom_array[10653] = 32'h00008949;
    // rom_array[10654] = 32'h00008951;
    // rom_array[10655] = 32'h00008959;
    // rom_array[10656] = 32'h00008961;
    // rom_array[10657] = 32'h00008969;
    // rom_array[10658] = 32'h00008971;
    // rom_array[10659] = 32'h00008979;
    // rom_array[10660] = 32'h00008981;
    // rom_array[10661] = 32'hFFFFFFF1;
    // rom_array[10662] = 32'hFFFFFFF1;
    // rom_array[10663] = 32'hFFFFFFF1;
    // rom_array[10664] = 32'hFFFFFFF1;
    // rom_array[10665] = 32'h00008989;
    // rom_array[10666] = 32'h00008991;
    // rom_array[10667] = 32'h00008999;
    // rom_array[10668] = 32'h000089a1;
    // rom_array[10669] = 32'h000089a9;
    // rom_array[10670] = 32'h000089b1;
    // rom_array[10671] = 32'h000089b9;
    // rom_array[10672] = 32'h000089c1;
    // rom_array[10673] = 32'hFFFFFFF0;
    // rom_array[10674] = 32'hFFFFFFF0;
    // rom_array[10675] = 32'hFFFFFFF0;
    // rom_array[10676] = 32'hFFFFFFF0;
    // rom_array[10677] = 32'h000089c9;
    // rom_array[10678] = 32'h000089d1;
    // rom_array[10679] = 32'hFFFFFFF0;
    // rom_array[10680] = 32'hFFFFFFF0;
    // rom_array[10681] = 32'h000089d9;
    // rom_array[10682] = 32'h000089e1;
    // rom_array[10683] = 32'h000089e9;
    // rom_array[10684] = 32'h000089f1;
    // rom_array[10685] = 32'h000089f9;
    // rom_array[10686] = 32'h00008a01;
    // rom_array[10687] = 32'h00008a09;
    // rom_array[10688] = 32'h00008a11;
    // rom_array[10689] = 32'h00008a19;
    // rom_array[10690] = 32'h00008a21;
    // rom_array[10691] = 32'hFFFFFFF0;
    // rom_array[10692] = 32'hFFFFFFF0;
    // rom_array[10693] = 32'h00008a29;
    // rom_array[10694] = 32'h00008a31;
    // rom_array[10695] = 32'hFFFFFFF0;
    // rom_array[10696] = 32'hFFFFFFF0;
    // rom_array[10697] = 32'h00008a39;
    // rom_array[10698] = 32'h00008a41;
    // rom_array[10699] = 32'h00008a49;
    // rom_array[10700] = 32'h00008a51;
    // rom_array[10701] = 32'hFFFFFFF1;
    // rom_array[10702] = 32'hFFFFFFF1;
    // rom_array[10703] = 32'hFFFFFFF1;
    // rom_array[10704] = 32'hFFFFFFF1;
    // rom_array[10705] = 32'h00008a59;
    // rom_array[10706] = 32'h00008a61;
    // rom_array[10707] = 32'h00008a69;
    // rom_array[10708] = 32'h00008a71;
    // rom_array[10709] = 32'hFFFFFFF1;
    // rom_array[10710] = 32'hFFFFFFF1;
    // rom_array[10711] = 32'hFFFFFFF1;
    // rom_array[10712] = 32'hFFFFFFF1;
    // rom_array[10713] = 32'h00008a79;
    // rom_array[10714] = 32'h00008a81;
    // rom_array[10715] = 32'hFFFFFFF1;
    // rom_array[10716] = 32'hFFFFFFF1;
    // rom_array[10717] = 32'h00008a89;
    // rom_array[10718] = 32'h00008a91;
    // rom_array[10719] = 32'hFFFFFFF1;
    // rom_array[10720] = 32'hFFFFFFF1;
    // rom_array[10721] = 32'h00008a99;
    // rom_array[10722] = 32'h00008aa1;
    // rom_array[10723] = 32'h00008aa9;
    // rom_array[10724] = 32'h00008ab1;
    // rom_array[10725] = 32'h00008ab9;
    // rom_array[10726] = 32'h00008ac1;
    // rom_array[10727] = 32'hFFFFFFF1;
    // rom_array[10728] = 32'hFFFFFFF1;
    // rom_array[10729] = 32'h00008ac9;
    // rom_array[10730] = 32'h00008ad1;
    // rom_array[10731] = 32'h00008ad9;
    // rom_array[10732] = 32'h00008ae1;
    // rom_array[10733] = 32'hFFFFFFF1;
    // rom_array[10734] = 32'hFFFFFFF1;
    // rom_array[10735] = 32'h00008ae9;
    // rom_array[10736] = 32'h00008af1;
    // rom_array[10737] = 32'h00008af9;
    // rom_array[10738] = 32'h00008b01;
    // rom_array[10739] = 32'hFFFFFFF1;
    // rom_array[10740] = 32'hFFFFFFF1;
    // rom_array[10741] = 32'h00008b09;
    // rom_array[10742] = 32'h00008b11;
    // rom_array[10743] = 32'hFFFFFFF1;
    // rom_array[10744] = 32'hFFFFFFF1;
    // rom_array[10745] = 32'hFFFFFFF1;
    // rom_array[10746] = 32'hFFFFFFF1;
    // rom_array[10747] = 32'h00008b19;
    // rom_array[10748] = 32'h00008b21;
    // rom_array[10749] = 32'hFFFFFFF1;
    // rom_array[10750] = 32'hFFFFFFF1;
    // rom_array[10751] = 32'h00008b29;
    // rom_array[10752] = 32'h00008b31;
    // rom_array[10753] = 32'h00008b39;
    // rom_array[10754] = 32'h00008b41;
    // rom_array[10755] = 32'h00008b49;
    // rom_array[10756] = 32'h00008b51;
    // rom_array[10757] = 32'hFFFFFFF0;
    // rom_array[10758] = 32'hFFFFFFF0;
    // rom_array[10759] = 32'hFFFFFFF0;
    // rom_array[10760] = 32'hFFFFFFF0;
    // rom_array[10761] = 32'h00008b59;
    // rom_array[10762] = 32'h00008b61;
    // rom_array[10763] = 32'h00008b69;
    // rom_array[10764] = 32'h00008b71;
    // rom_array[10765] = 32'hFFFFFFF1;
    // rom_array[10766] = 32'hFFFFFFF1;
    // rom_array[10767] = 32'h00008b79;
    // rom_array[10768] = 32'h00008b81;
    // rom_array[10769] = 32'h00008b89;
    // rom_array[10770] = 32'h00008b91;
    // rom_array[10771] = 32'h00008b99;
    // rom_array[10772] = 32'h00008ba1;
    // rom_array[10773] = 32'h00008ba9;
    // rom_array[10774] = 32'h00008bb1;
    // rom_array[10775] = 32'h00008bb9;
    // rom_array[10776] = 32'h00008bc1;
    // rom_array[10777] = 32'h00008bc9;
    // rom_array[10778] = 32'h00008bd1;
    // rom_array[10779] = 32'hFFFFFFF1;
    // rom_array[10780] = 32'hFFFFFFF1;
    // rom_array[10781] = 32'h00008bd9;
    // rom_array[10782] = 32'h00008be1;
    // rom_array[10783] = 32'h00008be9;
    // rom_array[10784] = 32'h00008bf1;
    // rom_array[10785] = 32'hFFFFFFF1;
    // rom_array[10786] = 32'hFFFFFFF1;
    // rom_array[10787] = 32'hFFFFFFF1;
    // rom_array[10788] = 32'hFFFFFFF1;
    // rom_array[10789] = 32'h00008bf9;
    // rom_array[10790] = 32'h00008c01;
    // rom_array[10791] = 32'h00008c09;
    // rom_array[10792] = 32'h00008c11;
    // rom_array[10793] = 32'hFFFFFFF1;
    // rom_array[10794] = 32'hFFFFFFF1;
    // rom_array[10795] = 32'hFFFFFFF1;
    // rom_array[10796] = 32'hFFFFFFF1;
    // rom_array[10797] = 32'h00008c19;
    // rom_array[10798] = 32'h00008c21;
    // rom_array[10799] = 32'h00008c29;
    // rom_array[10800] = 32'h00008c31;
    // rom_array[10801] = 32'hFFFFFFF1;
    // rom_array[10802] = 32'hFFFFFFF1;
    // rom_array[10803] = 32'hFFFFFFF1;
    // rom_array[10804] = 32'hFFFFFFF1;
    // rom_array[10805] = 32'h00008c39;
    // rom_array[10806] = 32'h00008c41;
    // rom_array[10807] = 32'h00008c49;
    // rom_array[10808] = 32'h00008c51;
    // rom_array[10809] = 32'hFFFFFFF1;
    // rom_array[10810] = 32'hFFFFFFF1;
    // rom_array[10811] = 32'h00008c59;
    // rom_array[10812] = 32'h00008c61;
    // rom_array[10813] = 32'h00008c69;
    // rom_array[10814] = 32'h00008c71;
    // rom_array[10815] = 32'h00008c79;
    // rom_array[10816] = 32'h00008c81;
    // rom_array[10817] = 32'hFFFFFFF0;
    // rom_array[10818] = 32'hFFFFFFF0;
    // rom_array[10819] = 32'hFFFFFFF0;
    // rom_array[10820] = 32'hFFFFFFF0;
    // rom_array[10821] = 32'h00008c89;
    // rom_array[10822] = 32'h00008c91;
    // rom_array[10823] = 32'h00008c99;
    // rom_array[10824] = 32'h00008ca1;
    // rom_array[10825] = 32'hFFFFFFF0;
    // rom_array[10826] = 32'hFFFFFFF0;
    // rom_array[10827] = 32'hFFFFFFF0;
    // rom_array[10828] = 32'hFFFFFFF0;
    // rom_array[10829] = 32'h00008ca9;
    // rom_array[10830] = 32'h00008cb1;
    // rom_array[10831] = 32'h00008cb9;
    // rom_array[10832] = 32'h00008cc1;
    // rom_array[10833] = 32'h00008cc9;
    // rom_array[10834] = 32'h00008cd1;
    // rom_array[10835] = 32'hFFFFFFF1;
    // rom_array[10836] = 32'hFFFFFFF1;
    // rom_array[10837] = 32'h00008cd9;
    // rom_array[10838] = 32'h00008ce1;
    // rom_array[10839] = 32'hFFFFFFF1;
    // rom_array[10840] = 32'hFFFFFFF1;
    // rom_array[10841] = 32'h00008ce9;
    // rom_array[10842] = 32'h00008cf1;
    // rom_array[10843] = 32'hFFFFFFF1;
    // rom_array[10844] = 32'hFFFFFFF1;
    // rom_array[10845] = 32'h00008cf9;
    // rom_array[10846] = 32'h00008d01;
    // rom_array[10847] = 32'hFFFFFFF1;
    // rom_array[10848] = 32'hFFFFFFF1;
    // rom_array[10849] = 32'h00008d09;
    // rom_array[10850] = 32'h00008d11;
    // rom_array[10851] = 32'hFFFFFFF1;
    // rom_array[10852] = 32'hFFFFFFF1;
    // rom_array[10853] = 32'h00008d19;
    // rom_array[10854] = 32'h00008d21;
    // rom_array[10855] = 32'hFFFFFFF1;
    // rom_array[10856] = 32'hFFFFFFF1;
    // rom_array[10857] = 32'hFFFFFFF0;
    // rom_array[10858] = 32'hFFFFFFF0;
    // rom_array[10859] = 32'hFFFFFFF0;
    // rom_array[10860] = 32'hFFFFFFF0;
    // rom_array[10861] = 32'h00008d29;
    // rom_array[10862] = 32'h00008d31;
    // rom_array[10863] = 32'hFFFFFFF0;
    // rom_array[10864] = 32'hFFFFFFF0;
    // rom_array[10865] = 32'h00008d39;
    // rom_array[10866] = 32'h00008d41;
    // rom_array[10867] = 32'hFFFFFFF0;
    // rom_array[10868] = 32'hFFFFFFF0;
    // rom_array[10869] = 32'h00008d49;
    // rom_array[10870] = 32'h00008d51;
    // rom_array[10871] = 32'hFFFFFFF0;
    // rom_array[10872] = 32'hFFFFFFF0;
    // rom_array[10873] = 32'h00008d59;
    // rom_array[10874] = 32'h00008d61;
    // rom_array[10875] = 32'hFFFFFFF0;
    // rom_array[10876] = 32'hFFFFFFF0;
    // rom_array[10877] = 32'h00008d69;
    // rom_array[10878] = 32'h00008d71;
    // rom_array[10879] = 32'hFFFFFFF0;
    // rom_array[10880] = 32'hFFFFFFF0;
    // rom_array[10881] = 32'h00008d79;
    // rom_array[10882] = 32'h00008d81;
    // rom_array[10883] = 32'h00008d89;
    // rom_array[10884] = 32'h00008d91;
    // rom_array[10885] = 32'h00008d99;
    // rom_array[10886] = 32'h00008da1;
    // rom_array[10887] = 32'hFFFFFFF1;
    // rom_array[10888] = 32'hFFFFFFF1;
    // rom_array[10889] = 32'h00008da9;
    // rom_array[10890] = 32'h00008db1;
    // rom_array[10891] = 32'h00008db9;
    // rom_array[10892] = 32'h00008dc1;
    // rom_array[10893] = 32'hFFFFFFF1;
    // rom_array[10894] = 32'hFFFFFFF1;
    // rom_array[10895] = 32'hFFFFFFF1;
    // rom_array[10896] = 32'hFFFFFFF1;
    // rom_array[10897] = 32'h00008dc9;
    // rom_array[10898] = 32'h00008dd1;
    // rom_array[10899] = 32'h00008dd9;
    // rom_array[10900] = 32'h00008de1;
    // rom_array[10901] = 32'hFFFFFFF1;
    // rom_array[10902] = 32'hFFFFFFF1;
    // rom_array[10903] = 32'hFFFFFFF1;
    // rom_array[10904] = 32'hFFFFFFF1;
    // rom_array[10905] = 32'h00008de9;
    // rom_array[10906] = 32'h00008df1;
    // rom_array[10907] = 32'h00008df9;
    // rom_array[10908] = 32'h00008e01;
    // rom_array[10909] = 32'hFFFFFFF1;
    // rom_array[10910] = 32'hFFFFFFF1;
    // rom_array[10911] = 32'hFFFFFFF1;
    // rom_array[10912] = 32'hFFFFFFF1;
    // rom_array[10913] = 32'h00008e09;
    // rom_array[10914] = 32'h00008e11;
    // rom_array[10915] = 32'hFFFFFFF1;
    // rom_array[10916] = 32'hFFFFFFF1;
    // rom_array[10917] = 32'h00008e19;
    // rom_array[10918] = 32'h00008e21;
    // rom_array[10919] = 32'hFFFFFFF1;
    // rom_array[10920] = 32'hFFFFFFF1;
    // rom_array[10921] = 32'h00008e29;
    // rom_array[10922] = 32'h00008e31;
    // rom_array[10923] = 32'hFFFFFFF1;
    // rom_array[10924] = 32'hFFFFFFF1;
    // rom_array[10925] = 32'h00008e39;
    // rom_array[10926] = 32'h00008e41;
    // rom_array[10927] = 32'hFFFFFFF1;
    // rom_array[10928] = 32'hFFFFFFF1;
    // rom_array[10929] = 32'h00008e49;
    // rom_array[10930] = 32'h00008e51;
    // rom_array[10931] = 32'hFFFFFFF1;
    // rom_array[10932] = 32'hFFFFFFF1;
    // rom_array[10933] = 32'h00008e59;
    // rom_array[10934] = 32'h00008e61;
    // rom_array[10935] = 32'hFFFFFFF1;
    // rom_array[10936] = 32'hFFFFFFF1;
    // rom_array[10937] = 32'h00008e69;
    // rom_array[10938] = 32'h00008e71;
    // rom_array[10939] = 32'hFFFFFFF1;
    // rom_array[10940] = 32'hFFFFFFF1;
    // rom_array[10941] = 32'h00008e79;
    // rom_array[10942] = 32'h00008e81;
    // rom_array[10943] = 32'h00008e89;
    // rom_array[10944] = 32'h00008e91;
    // rom_array[10945] = 32'hFFFFFFF1;
    // rom_array[10946] = 32'hFFFFFFF1;
    // rom_array[10947] = 32'hFFFFFFF1;
    // rom_array[10948] = 32'hFFFFFFF1;
    // rom_array[10949] = 32'h00008e99;
    // rom_array[10950] = 32'h00008ea1;
    // rom_array[10951] = 32'h00008ea9;
    // rom_array[10952] = 32'h00008eb1;
    // rom_array[10953] = 32'h00008eb9;
    // rom_array[10954] = 32'h00008ec1;
    // rom_array[10955] = 32'hFFFFFFF1;
    // rom_array[10956] = 32'hFFFFFFF1;
    // rom_array[10957] = 32'h00008ec9;
    // rom_array[10958] = 32'h00008ed1;
    // rom_array[10959] = 32'hFFFFFFF1;
    // rom_array[10960] = 32'hFFFFFFF1;
    // rom_array[10961] = 32'h00008ed9;
    // rom_array[10962] = 32'h00008ee1;
    // rom_array[10963] = 32'h00008ee9;
    // rom_array[10964] = 32'h00008ef1;
    // rom_array[10965] = 32'h00008ef9;
    // rom_array[10966] = 32'h00008f01;
    // rom_array[10967] = 32'hFFFFFFF0;
    // rom_array[10968] = 32'hFFFFFFF0;
    // rom_array[10969] = 32'h00008f09;
    // rom_array[10970] = 32'h00008f11;
    // rom_array[10971] = 32'h00008f19;
    // rom_array[10972] = 32'h00008f21;
    // rom_array[10973] = 32'hFFFFFFF0;
    // rom_array[10974] = 32'hFFFFFFF0;
    // rom_array[10975] = 32'hFFFFFFF0;
    // rom_array[10976] = 32'hFFFFFFF0;
    // rom_array[10977] = 32'h00008f29;
    // rom_array[10978] = 32'h00008f31;
    // rom_array[10979] = 32'h00008f39;
    // rom_array[10980] = 32'h00008f41;
    // rom_array[10981] = 32'hFFFFFFF0;
    // rom_array[10982] = 32'hFFFFFFF0;
    // rom_array[10983] = 32'hFFFFFFF0;
    // rom_array[10984] = 32'hFFFFFFF0;
    // rom_array[10985] = 32'h00008f49;
    // rom_array[10986] = 32'h00008f51;
    // rom_array[10987] = 32'h00008f59;
    // rom_array[10988] = 32'h00008f61;
    // rom_array[10989] = 32'hFFFFFFF0;
    // rom_array[10990] = 32'hFFFFFFF0;
    // rom_array[10991] = 32'hFFFFFFF0;
    // rom_array[10992] = 32'hFFFFFFF0;
    // rom_array[10993] = 32'h00008f69;
    // rom_array[10994] = 32'h00008f71;
    // rom_array[10995] = 32'hFFFFFFF0;
    // rom_array[10996] = 32'hFFFFFFF0;
    // rom_array[10997] = 32'h00008f79;
    // rom_array[10998] = 32'h00008f81;
    // rom_array[10999] = 32'hFFFFFFF0;
    // rom_array[11000] = 32'hFFFFFFF0;
    // rom_array[11001] = 32'h00008f89;
    // rom_array[11002] = 32'h00008f91;
    // rom_array[11003] = 32'hFFFFFFF0;
    // rom_array[11004] = 32'hFFFFFFF0;
    // rom_array[11005] = 32'h00008f99;
    // rom_array[11006] = 32'h00008fa1;
    // rom_array[11007] = 32'hFFFFFFF0;
    // rom_array[11008] = 32'hFFFFFFF0;
    // rom_array[11009] = 32'h00008fa9;
    // rom_array[11010] = 32'h00008fb1;
    // rom_array[11011] = 32'h00008fb9;
    // rom_array[11012] = 32'h00008fc1;
    // rom_array[11013] = 32'h00008fc9;
    // rom_array[11014] = 32'h00008fd1;
    // rom_array[11015] = 32'h00008fd9;
    // rom_array[11016] = 32'h00008fe1;
    // rom_array[11017] = 32'h00008fe9;
    // rom_array[11018] = 32'h00008ff1;
    // rom_array[11019] = 32'h00008ff9;
    // rom_array[11020] = 32'h00009001;
    // rom_array[11021] = 32'h00009009;
    // rom_array[11022] = 32'h00009011;
    // rom_array[11023] = 32'hFFFFFFF1;
    // rom_array[11024] = 32'hFFFFFFF1;
    // rom_array[11025] = 32'h00009019;
    // rom_array[11026] = 32'h00009021;
    // rom_array[11027] = 32'hFFFFFFF1;
    // rom_array[11028] = 32'hFFFFFFF1;
    // rom_array[11029] = 32'h00009029;
    // rom_array[11030] = 32'h00009031;
    // rom_array[11031] = 32'h00009039;
    // rom_array[11032] = 32'h00009041;
    // rom_array[11033] = 32'h00009049;
    // rom_array[11034] = 32'h00009051;
    // rom_array[11035] = 32'hFFFFFFF0;
    // rom_array[11036] = 32'hFFFFFFF0;
    // rom_array[11037] = 32'h00009059;
    // rom_array[11038] = 32'h00009061;
    // rom_array[11039] = 32'hFFFFFFF0;
    // rom_array[11040] = 32'hFFFFFFF0;
    // rom_array[11041] = 32'h00009069;
    // rom_array[11042] = 32'h00009071;
    // rom_array[11043] = 32'h00009079;
    // rom_array[11044] = 32'h00009081;
    // rom_array[11045] = 32'h00009089;
    // rom_array[11046] = 32'h00009091;
    // rom_array[11047] = 32'hFFFFFFF1;
    // rom_array[11048] = 32'hFFFFFFF1;
    // rom_array[11049] = 32'h00009099;
    // rom_array[11050] = 32'h000090a1;
    // rom_array[11051] = 32'hFFFFFFF0;
    // rom_array[11052] = 32'hFFFFFFF0;
    // rom_array[11053] = 32'hFFFFFFF0;
    // rom_array[11054] = 32'hFFFFFFF0;
    // rom_array[11055] = 32'hFFFFFFF0;
    // rom_array[11056] = 32'hFFFFFFF0;
    // rom_array[11057] = 32'h000090a9;
    // rom_array[11058] = 32'h000090b1;
    // rom_array[11059] = 32'hFFFFFFF1;
    // rom_array[11060] = 32'hFFFFFFF1;
    // rom_array[11061] = 32'h000090b9;
    // rom_array[11062] = 32'h000090c1;
    // rom_array[11063] = 32'hFFFFFFF1;
    // rom_array[11064] = 32'hFFFFFFF1;
    // rom_array[11065] = 32'h000090c9;
    // rom_array[11066] = 32'h000090d1;
    // rom_array[11067] = 32'h000090d9;
    // rom_array[11068] = 32'h000090e1;
    // rom_array[11069] = 32'hFFFFFFF1;
    // rom_array[11070] = 32'hFFFFFFF1;
    // rom_array[11071] = 32'hFFFFFFF1;
    // rom_array[11072] = 32'hFFFFFFF1;
    // rom_array[11073] = 32'h000090e9;
    // rom_array[11074] = 32'h000090f1;
    // rom_array[11075] = 32'h000090f9;
    // rom_array[11076] = 32'h00009101;
    // rom_array[11077] = 32'hFFFFFFF1;
    // rom_array[11078] = 32'hFFFFFFF1;
    // rom_array[11079] = 32'hFFFFFFF1;
    // rom_array[11080] = 32'hFFFFFFF1;
    // rom_array[11081] = 32'h00009109;
    // rom_array[11082] = 32'h00009111;
    // rom_array[11083] = 32'h00009119;
    // rom_array[11084] = 32'h00009121;
    // rom_array[11085] = 32'hFFFFFFF1;
    // rom_array[11086] = 32'hFFFFFFF1;
    // rom_array[11087] = 32'hFFFFFFF1;
    // rom_array[11088] = 32'hFFFFFFF1;
    // rom_array[11089] = 32'h00009129;
    // rom_array[11090] = 32'h00009131;
    // rom_array[11091] = 32'h00009139;
    // rom_array[11092] = 32'h00009141;
    // rom_array[11093] = 32'hFFFFFFF1;
    // rom_array[11094] = 32'hFFFFFFF1;
    // rom_array[11095] = 32'hFFFFFFF1;
    // rom_array[11096] = 32'hFFFFFFF1;
    // rom_array[11097] = 32'hFFFFFFF0;
    // rom_array[11098] = 32'hFFFFFFF0;
    // rom_array[11099] = 32'hFFFFFFF0;
    // rom_array[11100] = 32'hFFFFFFF0;
    // rom_array[11101] = 32'h00009149;
    // rom_array[11102] = 32'h00009151;
    // rom_array[11103] = 32'h00009159;
    // rom_array[11104] = 32'h00009161;
    // rom_array[11105] = 32'hFFFFFFF0;
    // rom_array[11106] = 32'hFFFFFFF0;
    // rom_array[11107] = 32'hFFFFFFF0;
    // rom_array[11108] = 32'hFFFFFFF0;
    // rom_array[11109] = 32'h00009169;
    // rom_array[11110] = 32'h00009171;
    // rom_array[11111] = 32'h00009179;
    // rom_array[11112] = 32'h00009181;
    // rom_array[11113] = 32'h00009189;
    // rom_array[11114] = 32'h00009191;
    // rom_array[11115] = 32'hFFFFFFF1;
    // rom_array[11116] = 32'hFFFFFFF1;
    // rom_array[11117] = 32'h00009199;
    // rom_array[11118] = 32'h000091a1;
    // rom_array[11119] = 32'hFFFFFFF1;
    // rom_array[11120] = 32'hFFFFFFF1;
    // rom_array[11121] = 32'hFFFFFFF0;
    // rom_array[11122] = 32'hFFFFFFF0;
    // rom_array[11123] = 32'hFFFFFFF0;
    // rom_array[11124] = 32'hFFFFFFF0;
    // rom_array[11125] = 32'h000091a9;
    // rom_array[11126] = 32'h000091b1;
    // rom_array[11127] = 32'hFFFFFFF0;
    // rom_array[11128] = 32'hFFFFFFF0;
    // rom_array[11129] = 32'h000091b9;
    // rom_array[11130] = 32'h000091c1;
    // rom_array[11131] = 32'hFFFFFFF0;
    // rom_array[11132] = 32'hFFFFFFF0;
    // rom_array[11133] = 32'h000091c9;
    // rom_array[11134] = 32'h000091d1;
    // rom_array[11135] = 32'hFFFFFFF0;
    // rom_array[11136] = 32'hFFFFFFF0;
    // rom_array[11137] = 32'h000091d9;
    // rom_array[11138] = 32'h000091e1;
    // rom_array[11139] = 32'h000091e9;
    // rom_array[11140] = 32'h000091f1;
    // rom_array[11141] = 32'h000091f9;
    // rom_array[11142] = 32'h00009201;
    // rom_array[11143] = 32'hFFFFFFF1;
    // rom_array[11144] = 32'hFFFFFFF1;
    // rom_array[11145] = 32'h00009209;
    // rom_array[11146] = 32'h00009211;
    // rom_array[11147] = 32'h00009219;
    // rom_array[11148] = 32'h00009221;
    // rom_array[11149] = 32'hFFFFFFF1;
    // rom_array[11150] = 32'hFFFFFFF1;
    // rom_array[11151] = 32'hFFFFFFF1;
    // rom_array[11152] = 32'hFFFFFFF1;
    // rom_array[11153] = 32'h00009229;
    // rom_array[11154] = 32'h00009231;
    // rom_array[11155] = 32'hFFFFFFF1;
    // rom_array[11156] = 32'hFFFFFFF1;
    // rom_array[11157] = 32'h00009239;
    // rom_array[11158] = 32'h00009241;
    // rom_array[11159] = 32'hFFFFFFF1;
    // rom_array[11160] = 32'hFFFFFFF1;
    // rom_array[11161] = 32'h00009249;
    // rom_array[11162] = 32'h00009251;
    // rom_array[11163] = 32'h00009259;
    // rom_array[11164] = 32'h00009261;
    // rom_array[11165] = 32'h00009269;
    // rom_array[11166] = 32'h00009271;
    // rom_array[11167] = 32'hFFFFFFF1;
    // rom_array[11168] = 32'hFFFFFFF1;
    // rom_array[11169] = 32'h00009279;
    // rom_array[11170] = 32'h00009281;
    // rom_array[11171] = 32'h00009289;
    // rom_array[11172] = 32'h00009291;
    // rom_array[11173] = 32'hFFFFFFF0;
    // rom_array[11174] = 32'hFFFFFFF0;
    // rom_array[11175] = 32'hFFFFFFF0;
    // rom_array[11176] = 32'hFFFFFFF0;
    // rom_array[11177] = 32'h00009299;
    // rom_array[11178] = 32'h000092a1;
    // rom_array[11179] = 32'hFFFFFFF1;
    // rom_array[11180] = 32'hFFFFFFF1;
    // rom_array[11181] = 32'h000092a9;
    // rom_array[11182] = 32'h000092b1;
    // rom_array[11183] = 32'hFFFFFFF1;
    // rom_array[11184] = 32'hFFFFFFF1;
    // rom_array[11185] = 32'h000092b9;
    // rom_array[11186] = 32'h000092c1;
    // rom_array[11187] = 32'h000092c9;
    // rom_array[11188] = 32'h000092d1;
    // rom_array[11189] = 32'h000092d9;
    // rom_array[11190] = 32'h000092e1;
    // rom_array[11191] = 32'hFFFFFFF1;
    // rom_array[11192] = 32'hFFFFFFF1;
    // rom_array[11193] = 32'h000092e9;
    // rom_array[11194] = 32'h000092f1;
    // rom_array[11195] = 32'h000092f9;
    // rom_array[11196] = 32'h00009301;
    // rom_array[11197] = 32'hFFFFFFF1;
    // rom_array[11198] = 32'hFFFFFFF1;
    // rom_array[11199] = 32'hFFFFFFF1;
    // rom_array[11200] = 32'hFFFFFFF1;
    // rom_array[11201] = 32'h00009309;
    // rom_array[11202] = 32'h00009311;
    // rom_array[11203] = 32'hFFFFFFF1;
    // rom_array[11204] = 32'hFFFFFFF1;
    // rom_array[11205] = 32'h00009319;
    // rom_array[11206] = 32'h00009321;
    // rom_array[11207] = 32'hFFFFFFF1;
    // rom_array[11208] = 32'hFFFFFFF1;
    // rom_array[11209] = 32'h00009329;
    // rom_array[11210] = 32'h00009331;
    // rom_array[11211] = 32'h00009339;
    // rom_array[11212] = 32'h00009341;
    // rom_array[11213] = 32'h00009349;
    // rom_array[11214] = 32'h00009351;
    // rom_array[11215] = 32'hFFFFFFF1;
    // rom_array[11216] = 32'hFFFFFFF1;
    // rom_array[11217] = 32'h00009359;
    // rom_array[11218] = 32'h00009361;
    // rom_array[11219] = 32'h00009369;
    // rom_array[11220] = 32'h00009371;
    // rom_array[11221] = 32'hFFFFFFF1;
    // rom_array[11222] = 32'hFFFFFFF1;
    // rom_array[11223] = 32'hFFFFFFF1;
    // rom_array[11224] = 32'hFFFFFFF1;
    // rom_array[11225] = 32'h00009379;
    // rom_array[11226] = 32'h00009381;
    // rom_array[11227] = 32'hFFFFFFF0;
    // rom_array[11228] = 32'hFFFFFFF0;
    // rom_array[11229] = 32'h00009389;
    // rom_array[11230] = 32'h00009391;
    // rom_array[11231] = 32'hFFFFFFF0;
    // rom_array[11232] = 32'hFFFFFFF0;
    // rom_array[11233] = 32'h00009399;
    // rom_array[11234] = 32'h000093a1;
    // rom_array[11235] = 32'h000093a9;
    // rom_array[11236] = 32'h000093b1;
    // rom_array[11237] = 32'h000093b9;
    // rom_array[11238] = 32'h000093c1;
    // rom_array[11239] = 32'hFFFFFFF1;
    // rom_array[11240] = 32'hFFFFFFF1;
    // rom_array[11241] = 32'h000093c9;
    // rom_array[11242] = 32'h000093d1;
    // rom_array[11243] = 32'h000093d9;
    // rom_array[11244] = 32'h000093e1;
    // rom_array[11245] = 32'hFFFFFFF0;
    // rom_array[11246] = 32'hFFFFFFF0;
    // rom_array[11247] = 32'hFFFFFFF0;
    // rom_array[11248] = 32'hFFFFFFF0;
    // rom_array[11249] = 32'h000093e9;
    // rom_array[11250] = 32'h000093f1;
    // rom_array[11251] = 32'hFFFFFFF1;
    // rom_array[11252] = 32'hFFFFFFF1;
    // rom_array[11253] = 32'h000093f9;
    // rom_array[11254] = 32'h00009401;
    // rom_array[11255] = 32'h00009409;
    // rom_array[11256] = 32'h00009411;
    // rom_array[11257] = 32'hFFFFFFF1;
    // rom_array[11258] = 32'hFFFFFFF1;
    // rom_array[11259] = 32'hFFFFFFF1;
    // rom_array[11260] = 32'hFFFFFFF1;
    // rom_array[11261] = 32'h00009419;
    // rom_array[11262] = 32'h00009421;
    // rom_array[11263] = 32'h00009429;
    // rom_array[11264] = 32'h00009431;
    // rom_array[11265] = 32'h00009439;
    // rom_array[11266] = 32'h00009441;
    // rom_array[11267] = 32'h00009449;
    // rom_array[11268] = 32'h00009451;
    // rom_array[11269] = 32'h00009459;
    // rom_array[11270] = 32'h00009461;
    // rom_array[11271] = 32'hFFFFFFF0;
    // rom_array[11272] = 32'hFFFFFFF0;
    // rom_array[11273] = 32'h00009469;
    // rom_array[11274] = 32'h00009471;
    // rom_array[11275] = 32'h00009479;
    // rom_array[11276] = 32'h00009481;
    // rom_array[11277] = 32'hFFFFFFF0;
    // rom_array[11278] = 32'hFFFFFFF0;
    // rom_array[11279] = 32'hFFFFFFF0;
    // rom_array[11280] = 32'hFFFFFFF0;
    // rom_array[11281] = 32'h00009489;
    // rom_array[11282] = 32'h00009491;
    // rom_array[11283] = 32'hFFFFFFF0;
    // rom_array[11284] = 32'hFFFFFFF0;
    // rom_array[11285] = 32'h00009499;
    // rom_array[11286] = 32'h000094a1;
    // rom_array[11287] = 32'hFFFFFFF0;
    // rom_array[11288] = 32'hFFFFFFF0;
    // rom_array[11289] = 32'h000094a9;
    // rom_array[11290] = 32'h000094b1;
    // rom_array[11291] = 32'h000094b9;
    // rom_array[11292] = 32'h000094c1;
    // rom_array[11293] = 32'h000094c9;
    // rom_array[11294] = 32'h000094d1;
    // rom_array[11295] = 32'h000094d9;
    // rom_array[11296] = 32'h000094e1;
    // rom_array[11297] = 32'h000094e9;
    // rom_array[11298] = 32'h000094f1;
    // rom_array[11299] = 32'hFFFFFFF0;
    // rom_array[11300] = 32'hFFFFFFF0;
    // rom_array[11301] = 32'h000094f9;
    // rom_array[11302] = 32'h00009501;
    // rom_array[11303] = 32'hFFFFFFF0;
    // rom_array[11304] = 32'hFFFFFFF0;
    // rom_array[11305] = 32'h00009509;
    // rom_array[11306] = 32'h00009511;
    // rom_array[11307] = 32'hFFFFFFF1;
    // rom_array[11308] = 32'hFFFFFFF1;
    // rom_array[11309] = 32'h00009519;
    // rom_array[11310] = 32'h00009521;
    // rom_array[11311] = 32'h00009529;
    // rom_array[11312] = 32'h00009531;
    // rom_array[11313] = 32'h00009539;
    // rom_array[11314] = 32'h00009541;
    // rom_array[11315] = 32'hFFFFFFF0;
    // rom_array[11316] = 32'hFFFFFFF0;
    // rom_array[11317] = 32'h00009549;
    // rom_array[11318] = 32'h00009551;
    // rom_array[11319] = 32'hFFFFFFF0;
    // rom_array[11320] = 32'hFFFFFFF0;
    // rom_array[11321] = 32'h00009559;
    // rom_array[11322] = 32'h00009561;
    // rom_array[11323] = 32'h00009569;
    // rom_array[11324] = 32'h00009571;
    // rom_array[11325] = 32'hFFFFFFF0;
    // rom_array[11326] = 32'hFFFFFFF0;
    // rom_array[11327] = 32'hFFFFFFF0;
    // rom_array[11328] = 32'hFFFFFFF0;
    // rom_array[11329] = 32'h00009579;
    // rom_array[11330] = 32'h00009581;
    // rom_array[11331] = 32'h00009589;
    // rom_array[11332] = 32'h00009591;
    // rom_array[11333] = 32'hFFFFFFF0;
    // rom_array[11334] = 32'hFFFFFFF0;
    // rom_array[11335] = 32'hFFFFFFF0;
    // rom_array[11336] = 32'hFFFFFFF0;
    // rom_array[11337] = 32'h00009599;
    // rom_array[11338] = 32'h000095a1;
    // rom_array[11339] = 32'h000095a9;
    // rom_array[11340] = 32'h000095b1;
    // rom_array[11341] = 32'hFFFFFFF0;
    // rom_array[11342] = 32'hFFFFFFF0;
    // rom_array[11343] = 32'hFFFFFFF0;
    // rom_array[11344] = 32'hFFFFFFF0;
    // rom_array[11345] = 32'h000095b9;
    // rom_array[11346] = 32'h000095c1;
    // rom_array[11347] = 32'h000095c9;
    // rom_array[11348] = 32'h000095d1;
    // rom_array[11349] = 32'hFFFFFFF0;
    // rom_array[11350] = 32'hFFFFFFF0;
    // rom_array[11351] = 32'hFFFFFFF0;
    // rom_array[11352] = 32'hFFFFFFF0;
    // rom_array[11353] = 32'h000095d9;
    // rom_array[11354] = 32'h000095e1;
    // rom_array[11355] = 32'h000095e9;
    // rom_array[11356] = 32'h000095f1;
    // rom_array[11357] = 32'hFFFFFFF0;
    // rom_array[11358] = 32'hFFFFFFF0;
    // rom_array[11359] = 32'hFFFFFFF0;
    // rom_array[11360] = 32'hFFFFFFF0;
    // rom_array[11361] = 32'h000095f9;
    // rom_array[11362] = 32'h00009601;
    // rom_array[11363] = 32'h00009609;
    // rom_array[11364] = 32'h00009611;
    // rom_array[11365] = 32'hFFFFFFF0;
    // rom_array[11366] = 32'hFFFFFFF0;
    // rom_array[11367] = 32'hFFFFFFF0;
    // rom_array[11368] = 32'hFFFFFFF0;
    // rom_array[11369] = 32'h00009619;
    // rom_array[11370] = 32'h00009621;
    // rom_array[11371] = 32'h00009629;
    // rom_array[11372] = 32'h00009631;
    // rom_array[11373] = 32'h00009639;
    // rom_array[11374] = 32'h00009641;
    // rom_array[11375] = 32'hFFFFFFF1;
    // rom_array[11376] = 32'hFFFFFFF1;
    // rom_array[11377] = 32'h00009649;
    // rom_array[11378] = 32'h00009651;
    // rom_array[11379] = 32'h00009659;
    // rom_array[11380] = 32'h00009661;
    // rom_array[11381] = 32'hFFFFFFF1;
    // rom_array[11382] = 32'hFFFFFFF1;
    // rom_array[11383] = 32'hFFFFFFF1;
    // rom_array[11384] = 32'hFFFFFFF1;
    // rom_array[11385] = 32'h00009669;
    // rom_array[11386] = 32'h00009671;
    // rom_array[11387] = 32'hFFFFFFF1;
    // rom_array[11388] = 32'hFFFFFFF1;
    // rom_array[11389] = 32'h00009679;
    // rom_array[11390] = 32'h00009681;
    // rom_array[11391] = 32'hFFFFFFF1;
    // rom_array[11392] = 32'hFFFFFFF1;
    // rom_array[11393] = 32'h00009689;
    // rom_array[11394] = 32'h00009691;
    // rom_array[11395] = 32'h00009699;
    // rom_array[11396] = 32'h000096a1;
    // rom_array[11397] = 32'hFFFFFFF1;
    // rom_array[11398] = 32'hFFFFFFF1;
    // rom_array[11399] = 32'hFFFFFFF1;
    // rom_array[11400] = 32'hFFFFFFF1;
    // rom_array[11401] = 32'h000096a9;
    // rom_array[11402] = 32'h000096b1;
    // rom_array[11403] = 32'h000096b9;
    // rom_array[11404] = 32'h000096c1;
    // rom_array[11405] = 32'hFFFFFFF1;
    // rom_array[11406] = 32'hFFFFFFF1;
    // rom_array[11407] = 32'hFFFFFFF1;
    // rom_array[11408] = 32'hFFFFFFF1;
    // rom_array[11409] = 32'h000096c9;
    // rom_array[11410] = 32'h000096d1;
    // rom_array[11411] = 32'h000096d9;
    // rom_array[11412] = 32'h000096e1;
    // rom_array[11413] = 32'hFFFFFFF1;
    // rom_array[11414] = 32'hFFFFFFF1;
    // rom_array[11415] = 32'hFFFFFFF1;
    // rom_array[11416] = 32'hFFFFFFF1;
    // rom_array[11417] = 32'h000096e9;
    // rom_array[11418] = 32'h000096f1;
    // rom_array[11419] = 32'h000096f9;
    // rom_array[11420] = 32'h00009701;
    // rom_array[11421] = 32'hFFFFFFF1;
    // rom_array[11422] = 32'hFFFFFFF1;
    // rom_array[11423] = 32'hFFFFFFF1;
    // rom_array[11424] = 32'hFFFFFFF1;
    // rom_array[11425] = 32'h00009709;
    // rom_array[11426] = 32'h00009711;
    // rom_array[11427] = 32'h00009719;
    // rom_array[11428] = 32'h00009721;
    // rom_array[11429] = 32'h00009729;
    // rom_array[11430] = 32'h00009731;
    // rom_array[11431] = 32'hFFFFFFF1;
    // rom_array[11432] = 32'hFFFFFFF1;
    // rom_array[11433] = 32'h00009739;
    // rom_array[11434] = 32'h00009741;
    // rom_array[11435] = 32'h00009749;
    // rom_array[11436] = 32'h00009751;
    // rom_array[11437] = 32'hFFFFFFF1;
    // rom_array[11438] = 32'hFFFFFFF1;
    // rom_array[11439] = 32'hFFFFFFF1;
    // rom_array[11440] = 32'hFFFFFFF1;
    // rom_array[11441] = 32'h00009759;
    // rom_array[11442] = 32'h00009761;
    // rom_array[11443] = 32'hFFFFFFF1;
    // rom_array[11444] = 32'hFFFFFFF1;
    // rom_array[11445] = 32'h00009769;
    // rom_array[11446] = 32'h00009771;
    // rom_array[11447] = 32'hFFFFFFF1;
    // rom_array[11448] = 32'hFFFFFFF1;
    // rom_array[11449] = 32'h00009779;
    // rom_array[11450] = 32'h00009781;
    // rom_array[11451] = 32'hFFFFFFF1;
    // rom_array[11452] = 32'hFFFFFFF1;
    // rom_array[11453] = 32'h00009789;
    // rom_array[11454] = 32'h00009791;
    // rom_array[11455] = 32'hFFFFFFF1;
    // rom_array[11456] = 32'hFFFFFFF1;
    // rom_array[11457] = 32'h00009799;
    // rom_array[11458] = 32'h000097a1;
    // rom_array[11459] = 32'hFFFFFFF1;
    // rom_array[11460] = 32'hFFFFFFF1;
    // rom_array[11461] = 32'h000097a9;
    // rom_array[11462] = 32'h000097b1;
    // rom_array[11463] = 32'hFFFFFFF1;
    // rom_array[11464] = 32'hFFFFFFF1;
    // rom_array[11465] = 32'h000097b9;
    // rom_array[11466] = 32'h000097c1;
    // rom_array[11467] = 32'h000097c9;
    // rom_array[11468] = 32'h000097d1;
    // rom_array[11469] = 32'h000097d9;
    // rom_array[11470] = 32'h000097e1;
    // rom_array[11471] = 32'hFFFFFFF0;
    // rom_array[11472] = 32'hFFFFFFF0;
    // rom_array[11473] = 32'h000097e9;
    // rom_array[11474] = 32'h000097f1;
    // rom_array[11475] = 32'h000097f9;
    // rom_array[11476] = 32'h00009801;
    // rom_array[11477] = 32'hFFFFFFF0;
    // rom_array[11478] = 32'hFFFFFFF0;
    // rom_array[11479] = 32'hFFFFFFF0;
    // rom_array[11480] = 32'hFFFFFFF0;
    // rom_array[11481] = 32'h00009809;
    // rom_array[11482] = 32'h00009811;
    // rom_array[11483] = 32'hFFFFFFF0;
    // rom_array[11484] = 32'hFFFFFFF0;
    // rom_array[11485] = 32'h00009819;
    // rom_array[11486] = 32'h00009821;
    // rom_array[11487] = 32'hFFFFFFF0;
    // rom_array[11488] = 32'hFFFFFFF0;
    // rom_array[11489] = 32'h00009829;
    // rom_array[11490] = 32'h00009831;
    // rom_array[11491] = 32'h00009839;
    // rom_array[11492] = 32'h00009841;
    // rom_array[11493] = 32'hFFFFFFF0;
    // rom_array[11494] = 32'hFFFFFFF0;
    // rom_array[11495] = 32'hFFFFFFF0;
    // rom_array[11496] = 32'hFFFFFFF0;
    // rom_array[11497] = 32'h00009849;
    // rom_array[11498] = 32'h00009851;
    // rom_array[11499] = 32'h00009859;
    // rom_array[11500] = 32'h00009861;
    // rom_array[11501] = 32'hFFFFFFF0;
    // rom_array[11502] = 32'hFFFFFFF0;
    // rom_array[11503] = 32'hFFFFFFF0;
    // rom_array[11504] = 32'hFFFFFFF0;
    // rom_array[11505] = 32'h00009869;
    // rom_array[11506] = 32'h00009871;
    // rom_array[11507] = 32'hFFFFFFF0;
    // rom_array[11508] = 32'hFFFFFFF0;
    // rom_array[11509] = 32'h00009879;
    // rom_array[11510] = 32'h00009881;
    // rom_array[11511] = 32'hFFFFFFF0;
    // rom_array[11512] = 32'hFFFFFFF0;
    // rom_array[11513] = 32'h00009889;
    // rom_array[11514] = 32'h00009891;
    // rom_array[11515] = 32'hFFFFFFF0;
    // rom_array[11516] = 32'hFFFFFFF0;
    // rom_array[11517] = 32'h00009899;
    // rom_array[11518] = 32'h000098a1;
    // rom_array[11519] = 32'hFFFFFFF0;
    // rom_array[11520] = 32'hFFFFFFF0;
    // rom_array[11521] = 32'h000098a9;
    // rom_array[11522] = 32'h000098b1;
    // rom_array[11523] = 32'hFFFFFFF1;
    // rom_array[11524] = 32'hFFFFFFF1;
    // rom_array[11525] = 32'h000098b9;
    // rom_array[11526] = 32'h000098c1;
    // rom_array[11527] = 32'hFFFFFFF1;
    // rom_array[11528] = 32'hFFFFFFF1;
    // rom_array[11529] = 32'h000098c9;
    // rom_array[11530] = 32'h000098d1;
    // rom_array[11531] = 32'h000098d9;
    // rom_array[11532] = 32'h000098e1;
    // rom_array[11533] = 32'hFFFFFFF0;
    // rom_array[11534] = 32'hFFFFFFF0;
    // rom_array[11535] = 32'hFFFFFFF0;
    // rom_array[11536] = 32'hFFFFFFF0;
    // rom_array[11537] = 32'h000098e9;
    // rom_array[11538] = 32'h000098f1;
    // rom_array[11539] = 32'h000098f9;
    // rom_array[11540] = 32'h00009901;
    // rom_array[11541] = 32'hFFFFFFF0;
    // rom_array[11542] = 32'hFFFFFFF0;
    // rom_array[11543] = 32'hFFFFFFF0;
    // rom_array[11544] = 32'hFFFFFFF0;
    // rom_array[11545] = 32'h00009909;
    // rom_array[11546] = 32'h00009911;
    // rom_array[11547] = 32'hFFFFFFF0;
    // rom_array[11548] = 32'hFFFFFFF0;
    // rom_array[11549] = 32'h00009919;
    // rom_array[11550] = 32'h00009921;
    // rom_array[11551] = 32'hFFFFFFF0;
    // rom_array[11552] = 32'hFFFFFFF0;
    // rom_array[11553] = 32'h00009929;
    // rom_array[11554] = 32'h00009931;
    // rom_array[11555] = 32'hFFFFFFF0;
    // rom_array[11556] = 32'hFFFFFFF0;
    // rom_array[11557] = 32'hFFFFFFF0;
    // rom_array[11558] = 32'hFFFFFFF0;
    // rom_array[11559] = 32'hFFFFFFF0;
    // rom_array[11560] = 32'hFFFFFFF0;
    // rom_array[11561] = 32'h00009939;
    // rom_array[11562] = 32'h00009941;
    // rom_array[11563] = 32'h00009949;
    // rom_array[11564] = 32'h00009951;
    // rom_array[11565] = 32'hFFFFFFF0;
    // rom_array[11566] = 32'hFFFFFFF0;
    // rom_array[11567] = 32'hFFFFFFF0;
    // rom_array[11568] = 32'hFFFFFFF0;
    // rom_array[11569] = 32'h00009959;
    // rom_array[11570] = 32'h00009961;
    // rom_array[11571] = 32'h00009969;
    // rom_array[11572] = 32'h00009971;
    // rom_array[11573] = 32'hFFFFFFF0;
    // rom_array[11574] = 32'hFFFFFFF0;
    // rom_array[11575] = 32'hFFFFFFF0;
    // rom_array[11576] = 32'hFFFFFFF0;
    // rom_array[11577] = 32'h00009979;
    // rom_array[11578] = 32'h00009981;
    // rom_array[11579] = 32'h00009989;
    // rom_array[11580] = 32'h00009991;
    // rom_array[11581] = 32'hFFFFFFF0;
    // rom_array[11582] = 32'hFFFFFFF0;
    // rom_array[11583] = 32'hFFFFFFF0;
    // rom_array[11584] = 32'hFFFFFFF0;
    // rom_array[11585] = 32'h00009999;
    // rom_array[11586] = 32'h000099a1;
    // rom_array[11587] = 32'hFFFFFFF0;
    // rom_array[11588] = 32'hFFFFFFF0;
    // rom_array[11589] = 32'hFFFFFFF0;
    // rom_array[11590] = 32'hFFFFFFF0;
    // rom_array[11591] = 32'hFFFFFFF0;
    // rom_array[11592] = 32'hFFFFFFF0;
    // rom_array[11593] = 32'h000099a9;
    // rom_array[11594] = 32'h000099b1;
    // rom_array[11595] = 32'h000099b9;
    // rom_array[11596] = 32'h000099c1;
    // rom_array[11597] = 32'hFFFFFFF1;
    // rom_array[11598] = 32'hFFFFFFF1;
    // rom_array[11599] = 32'hFFFFFFF1;
    // rom_array[11600] = 32'hFFFFFFF1;
    // rom_array[11601] = 32'h000099c9;
    // rom_array[11602] = 32'h000099d1;
    // rom_array[11603] = 32'h000099d9;
    // rom_array[11604] = 32'h000099e1;
    // rom_array[11605] = 32'hFFFFFFF1;
    // rom_array[11606] = 32'hFFFFFFF1;
    // rom_array[11607] = 32'hFFFFFFF1;
    // rom_array[11608] = 32'hFFFFFFF1;
    // rom_array[11609] = 32'h000099e9;
    // rom_array[11610] = 32'h000099f1;
    // rom_array[11611] = 32'h000099f9;
    // rom_array[11612] = 32'h00009a01;
    // rom_array[11613] = 32'hFFFFFFF1;
    // rom_array[11614] = 32'hFFFFFFF1;
    // rom_array[11615] = 32'hFFFFFFF1;
    // rom_array[11616] = 32'hFFFFFFF1;
    // rom_array[11617] = 32'h00009a09;
    // rom_array[11618] = 32'h00009a11;
    // rom_array[11619] = 32'h00009a19;
    // rom_array[11620] = 32'h00009a21;
    // rom_array[11621] = 32'hFFFFFFF1;
    // rom_array[11622] = 32'hFFFFFFF1;
    // rom_array[11623] = 32'hFFFFFFF1;
    // rom_array[11624] = 32'hFFFFFFF1;
    // rom_array[11625] = 32'h00009a29;
    // rom_array[11626] = 32'h00009a31;
    // rom_array[11627] = 32'h00009a39;
    // rom_array[11628] = 32'h00009a41;
    // rom_array[11629] = 32'h00009a49;
    // rom_array[11630] = 32'h00009a51;
    // rom_array[11631] = 32'hFFFFFFF0;
    // rom_array[11632] = 32'hFFFFFFF0;
    // rom_array[11633] = 32'h00009a59;
    // rom_array[11634] = 32'h00009a61;
    // rom_array[11635] = 32'h00009a69;
    // rom_array[11636] = 32'h00009a71;
    // rom_array[11637] = 32'hFFFFFFF0;
    // rom_array[11638] = 32'hFFFFFFF0;
    // rom_array[11639] = 32'hFFFFFFF0;
    // rom_array[11640] = 32'hFFFFFFF0;
    // rom_array[11641] = 32'h00009a79;
    // rom_array[11642] = 32'h00009a81;
    // rom_array[11643] = 32'h00009a89;
    // rom_array[11644] = 32'h00009a91;
    // rom_array[11645] = 32'hFFFFFFF0;
    // rom_array[11646] = 32'hFFFFFFF0;
    // rom_array[11647] = 32'hFFFFFFF0;
    // rom_array[11648] = 32'hFFFFFFF0;
    // rom_array[11649] = 32'h00009a99;
    // rom_array[11650] = 32'h00009aa1;
    // rom_array[11651] = 32'h00009aa9;
    // rom_array[11652] = 32'h00009ab1;
    // rom_array[11653] = 32'h00009ab9;
    // rom_array[11654] = 32'h00009ac1;
    // rom_array[11655] = 32'hFFFFFFF1;
    // rom_array[11656] = 32'hFFFFFFF1;
    // rom_array[11657] = 32'h00009ac9;
    // rom_array[11658] = 32'h00009ad1;
    // rom_array[11659] = 32'h00009ad9;
    // rom_array[11660] = 32'h00009ae1;
    // rom_array[11661] = 32'hFFFFFFF1;
    // rom_array[11662] = 32'hFFFFFFF1;
    // rom_array[11663] = 32'hFFFFFFF1;
    // rom_array[11664] = 32'hFFFFFFF1;
    // rom_array[11665] = 32'h00009ae9;
    // rom_array[11666] = 32'h00009af1;
    // rom_array[11667] = 32'hFFFFFFF0;
    // rom_array[11668] = 32'hFFFFFFF0;
    // rom_array[11669] = 32'h00009af9;
    // rom_array[11670] = 32'h00009b01;
    // rom_array[11671] = 32'hFFFFFFF0;
    // rom_array[11672] = 32'hFFFFFFF0;
    // rom_array[11673] = 32'h00009b09;
    // rom_array[11674] = 32'h00009b11;
    // rom_array[11675] = 32'hFFFFFFF0;
    // rom_array[11676] = 32'hFFFFFFF0;
    // rom_array[11677] = 32'h00009b19;
    // rom_array[11678] = 32'h00009b21;
    // rom_array[11679] = 32'hFFFFFFF0;
    // rom_array[11680] = 32'hFFFFFFF0;
    // rom_array[11681] = 32'h00009b29;
    // rom_array[11682] = 32'h00009b31;
    // rom_array[11683] = 32'h00009b39;
    // rom_array[11684] = 32'h00009b41;
    // rom_array[11685] = 32'hFFFFFFF1;
    // rom_array[11686] = 32'hFFFFFFF1;
    // rom_array[11687] = 32'hFFFFFFF1;
    // rom_array[11688] = 32'hFFFFFFF1;
    // rom_array[11689] = 32'h00009b49;
    // rom_array[11690] = 32'h00009b51;
    // rom_array[11691] = 32'hFFFFFFF0;
    // rom_array[11692] = 32'hFFFFFFF0;
    // rom_array[11693] = 32'h00009b59;
    // rom_array[11694] = 32'h00009b61;
    // rom_array[11695] = 32'hFFFFFFF0;
    // rom_array[11696] = 32'hFFFFFFF0;
    // rom_array[11697] = 32'h00009b69;
    // rom_array[11698] = 32'h00009b71;
    // rom_array[11699] = 32'hFFFFFFF0;
    // rom_array[11700] = 32'hFFFFFFF0;
    // rom_array[11701] = 32'h00009b79;
    // rom_array[11702] = 32'h00009b81;
    // rom_array[11703] = 32'hFFFFFFF0;
    // rom_array[11704] = 32'hFFFFFFF0;
    // rom_array[11705] = 32'h00009b89;
    // rom_array[11706] = 32'h00009b91;
    // rom_array[11707] = 32'hFFFFFFF0;
    // rom_array[11708] = 32'hFFFFFFF0;
    // rom_array[11709] = 32'h00009b99;
    // rom_array[11710] = 32'h00009ba1;
    // rom_array[11711] = 32'hFFFFFFF0;
    // rom_array[11712] = 32'hFFFFFFF0;
    // rom_array[11713] = 32'h00009ba9;
    // rom_array[11714] = 32'h00009bb1;
    // rom_array[11715] = 32'hFFFFFFF1;
    // rom_array[11716] = 32'hFFFFFFF1;
    // rom_array[11717] = 32'h00009bb9;
    // rom_array[11718] = 32'h00009bc1;
    // rom_array[11719] = 32'hFFFFFFF1;
    // rom_array[11720] = 32'hFFFFFFF1;
    // rom_array[11721] = 32'h00009bc9;
    // rom_array[11722] = 32'h00009bd1;
    // rom_array[11723] = 32'hFFFFFFF1;
    // rom_array[11724] = 32'hFFFFFFF1;
    // rom_array[11725] = 32'h00009bd9;
    // rom_array[11726] = 32'h00009be1;
    // rom_array[11727] = 32'hFFFFFFF1;
    // rom_array[11728] = 32'hFFFFFFF1;
    // rom_array[11729] = 32'h00009be9;
    // rom_array[11730] = 32'h00009bf1;
    // rom_array[11731] = 32'hFFFFFFF0;
    // rom_array[11732] = 32'hFFFFFFF0;
    // rom_array[11733] = 32'h00009bf9;
    // rom_array[11734] = 32'h00009c01;
    // rom_array[11735] = 32'h00009c09;
    // rom_array[11736] = 32'h00009c11;
    // rom_array[11737] = 32'hFFFFFFF0;
    // rom_array[11738] = 32'hFFFFFFF0;
    // rom_array[11739] = 32'hFFFFFFF0;
    // rom_array[11740] = 32'hFFFFFFF0;
    // rom_array[11741] = 32'h00009c19;
    // rom_array[11742] = 32'h00009c21;
    // rom_array[11743] = 32'h00009c29;
    // rom_array[11744] = 32'h00009c31;
    // rom_array[11745] = 32'h00009c39;
    // rom_array[11746] = 32'h00009c41;
    // rom_array[11747] = 32'hFFFFFFF0;
    // rom_array[11748] = 32'hFFFFFFF0;
    // rom_array[11749] = 32'hFFFFFFF0;
    // rom_array[11750] = 32'hFFFFFFF0;
    // rom_array[11751] = 32'hFFFFFFF0;
    // rom_array[11752] = 32'hFFFFFFF0;
    // rom_array[11753] = 32'hFFFFFFF0;
    // rom_array[11754] = 32'hFFFFFFF0;
    // rom_array[11755] = 32'hFFFFFFF0;
    // rom_array[11756] = 32'hFFFFFFF0;
    // rom_array[11757] = 32'h00009c49;
    // rom_array[11758] = 32'h00009c51;
    // rom_array[11759] = 32'h00009c59;
    // rom_array[11760] = 32'h00009c61;
    // rom_array[11761] = 32'h00009c69;
    // rom_array[11762] = 32'h00009c71;
    // rom_array[11763] = 32'hFFFFFFF1;
    // rom_array[11764] = 32'hFFFFFFF1;
    // rom_array[11765] = 32'h00009c79;
    // rom_array[11766] = 32'h00009c81;
    // rom_array[11767] = 32'h00009c89;
    // rom_array[11768] = 32'h00009c91;
    // rom_array[11769] = 32'h00009c99;
    // rom_array[11770] = 32'h00009ca1;
    // rom_array[11771] = 32'h00009ca9;
    // rom_array[11772] = 32'h00009cb1;
    // rom_array[11773] = 32'hFFFFFFF1;
    // rom_array[11774] = 32'hFFFFFFF1;
    // rom_array[11775] = 32'h00009cb9;
    // rom_array[11776] = 32'h00009cc1;
    // rom_array[11777] = 32'h00009cc9;
    // rom_array[11778] = 32'h00009cd1;
    // rom_array[11779] = 32'hFFFFFFF0;
    // rom_array[11780] = 32'hFFFFFFF0;
    // rom_array[11781] = 32'h00009cd9;
    // rom_array[11782] = 32'h00009ce1;
    // rom_array[11783] = 32'hFFFFFFF0;
    // rom_array[11784] = 32'hFFFFFFF0;
    // rom_array[11785] = 32'h00009ce9;
    // rom_array[11786] = 32'h00009cf1;
    // rom_array[11787] = 32'hFFFFFFF0;
    // rom_array[11788] = 32'hFFFFFFF0;
    // rom_array[11789] = 32'h00009cf9;
    // rom_array[11790] = 32'h00009d01;
    // rom_array[11791] = 32'hFFFFFFF0;
    // rom_array[11792] = 32'hFFFFFFF0;
    // rom_array[11793] = 32'h00009d09;
    // rom_array[11794] = 32'h00009d11;
    // rom_array[11795] = 32'hFFFFFFF0;
    // rom_array[11796] = 32'hFFFFFFF0;
    // rom_array[11797] = 32'h00009d19;
    // rom_array[11798] = 32'h00009d21;
    // rom_array[11799] = 32'hFFFFFFF0;
    // rom_array[11800] = 32'hFFFFFFF0;
    // rom_array[11801] = 32'h00009d29;
    // rom_array[11802] = 32'h00009d31;
    // rom_array[11803] = 32'h00009d39;
    // rom_array[11804] = 32'h00009d41;
    // rom_array[11805] = 32'hFFFFFFF0;
    // rom_array[11806] = 32'hFFFFFFF0;
    // rom_array[11807] = 32'hFFFFFFF0;
    // rom_array[11808] = 32'hFFFFFFF0;
    // rom_array[11809] = 32'h00009d49;
    // rom_array[11810] = 32'h00009d51;
    // rom_array[11811] = 32'hFFFFFFF0;
    // rom_array[11812] = 32'hFFFFFFF0;
    // rom_array[11813] = 32'hFFFFFFF0;
    // rom_array[11814] = 32'hFFFFFFF0;
    // rom_array[11815] = 32'hFFFFFFF0;
    // rom_array[11816] = 32'hFFFFFFF0;
    // rom_array[11817] = 32'hFFFFFFF1;
    // rom_array[11818] = 32'hFFFFFFF1;
    // rom_array[11819] = 32'hFFFFFFF1;
    // rom_array[11820] = 32'hFFFFFFF1;
    // rom_array[11821] = 32'h00009d59;
    // rom_array[11822] = 32'h00009d61;
    // rom_array[11823] = 32'h00009d69;
    // rom_array[11824] = 32'h00009d71;
    // rom_array[11825] = 32'hFFFFFFF1;
    // rom_array[11826] = 32'hFFFFFFF1;
    // rom_array[11827] = 32'hFFFFFFF1;
    // rom_array[11828] = 32'hFFFFFFF1;
    // rom_array[11829] = 32'h00009d79;
    // rom_array[11830] = 32'h00009d81;
    // rom_array[11831] = 32'h00009d89;
    // rom_array[11832] = 32'h00009d91;
    // rom_array[11833] = 32'hFFFFFFF1;
    // rom_array[11834] = 32'hFFFFFFF1;
    // rom_array[11835] = 32'hFFFFFFF1;
    // rom_array[11836] = 32'hFFFFFFF1;
    // rom_array[11837] = 32'h00009d99;
    // rom_array[11838] = 32'h00009da1;
    // rom_array[11839] = 32'h00009da9;
    // rom_array[11840] = 32'h00009db1;
    // rom_array[11841] = 32'hFFFFFFF1;
    // rom_array[11842] = 32'hFFFFFFF1;
    // rom_array[11843] = 32'h00009db9;
    // rom_array[11844] = 32'h00009dc1;
    // rom_array[11845] = 32'h00009dc9;
    // rom_array[11846] = 32'h00009dd1;
    // rom_array[11847] = 32'h00009dd9;
    // rom_array[11848] = 32'h00009de1;
    // rom_array[11849] = 32'hFFFFFFF0;
    // rom_array[11850] = 32'hFFFFFFF0;
    // rom_array[11851] = 32'hFFFFFFF0;
    // rom_array[11852] = 32'hFFFFFFF0;
    // rom_array[11853] = 32'h00009de9;
    // rom_array[11854] = 32'h00009df1;
    // rom_array[11855] = 32'h00009df9;
    // rom_array[11856] = 32'h00009e01;
    // rom_array[11857] = 32'h00009e09;
    // rom_array[11858] = 32'h00009e11;
    // rom_array[11859] = 32'hFFFFFFF1;
    // rom_array[11860] = 32'hFFFFFFF1;
    // rom_array[11861] = 32'h00009e19;
    // rom_array[11862] = 32'h00009e21;
    // rom_array[11863] = 32'hFFFFFFF1;
    // rom_array[11864] = 32'hFFFFFFF1;
    // rom_array[11865] = 32'h00009e29;
    // rom_array[11866] = 32'h00009e31;
    // rom_array[11867] = 32'h00009e39;
    // rom_array[11868] = 32'h00009e41;
    // rom_array[11869] = 32'hFFFFFFF1;
    // rom_array[11870] = 32'hFFFFFFF1;
    // rom_array[11871] = 32'hFFFFFFF1;
    // rom_array[11872] = 32'hFFFFFFF1;
    // rom_array[11873] = 32'h00009e49;
    // rom_array[11874] = 32'h00009e51;
    // rom_array[11875] = 32'h00009e59;
    // rom_array[11876] = 32'h00009e61;
    // rom_array[11877] = 32'hFFFFFFF1;
    // rom_array[11878] = 32'hFFFFFFF1;
    // rom_array[11879] = 32'hFFFFFFF1;
    // rom_array[11880] = 32'hFFFFFFF1;
    // rom_array[11881] = 32'h00009e69;
    // rom_array[11882] = 32'h00009e71;
    // rom_array[11883] = 32'hFFFFFFF1;
    // rom_array[11884] = 32'hFFFFFFF1;
    // rom_array[11885] = 32'h00009e79;
    // rom_array[11886] = 32'h00009e81;
    // rom_array[11887] = 32'hFFFFFFF1;
    // rom_array[11888] = 32'hFFFFFFF1;
    // rom_array[11889] = 32'h00009e89;
    // rom_array[11890] = 32'h00009e91;
    // rom_array[11891] = 32'h00009e99;
    // rom_array[11892] = 32'h00009ea1;
    // rom_array[11893] = 32'hFFFFFFF1;
    // rom_array[11894] = 32'hFFFFFFF1;
    // rom_array[11895] = 32'hFFFFFFF1;
    // rom_array[11896] = 32'hFFFFFFF1;
    // rom_array[11897] = 32'h00009ea9;
    // rom_array[11898] = 32'h00009eb1;
    // rom_array[11899] = 32'hFFFFFFF1;
    // rom_array[11900] = 32'hFFFFFFF1;
    // rom_array[11901] = 32'h00009eb9;
    // rom_array[11902] = 32'h00009ec1;
    // rom_array[11903] = 32'hFFFFFFF1;
    // rom_array[11904] = 32'hFFFFFFF1;
    // rom_array[11905] = 32'hFFFFFFF0;
    // rom_array[11906] = 32'hFFFFFFF0;
    // rom_array[11907] = 32'hFFFFFFF0;
    // rom_array[11908] = 32'hFFFFFFF0;
    // rom_array[11909] = 32'h00009ec9;
    // rom_array[11910] = 32'h00009ed1;
    // rom_array[11911] = 32'h00009ed9;
    // rom_array[11912] = 32'h00009ee1;
    // rom_array[11913] = 32'hFFFFFFF0;
    // rom_array[11914] = 32'hFFFFFFF0;
    // rom_array[11915] = 32'hFFFFFFF0;
    // rom_array[11916] = 32'hFFFFFFF0;
    // rom_array[11917] = 32'h00009ee9;
    // rom_array[11918] = 32'h00009ef1;
    // rom_array[11919] = 32'hFFFFFFF0;
    // rom_array[11920] = 32'hFFFFFFF0;
    // rom_array[11921] = 32'h00009ef9;
    // rom_array[11922] = 32'h00009f01;
    // rom_array[11923] = 32'hFFFFFFF0;
    // rom_array[11924] = 32'hFFFFFFF0;
    // rom_array[11925] = 32'h00009f09;
    // rom_array[11926] = 32'h00009f11;
    // rom_array[11927] = 32'hFFFFFFF0;
    // rom_array[11928] = 32'hFFFFFFF0;
    // rom_array[11929] = 32'h00009f19;
    // rom_array[11930] = 32'h00009f21;
    // rom_array[11931] = 32'hFFFFFFF0;
    // rom_array[11932] = 32'hFFFFFFF0;
    // rom_array[11933] = 32'h00009f29;
    // rom_array[11934] = 32'h00009f31;
    // rom_array[11935] = 32'hFFFFFFF0;
    // rom_array[11936] = 32'hFFFFFFF0;
    // rom_array[11937] = 32'h00009f39;
    // rom_array[11938] = 32'h00009f41;
    // rom_array[11939] = 32'hFFFFFFF0;
    // rom_array[11940] = 32'hFFFFFFF0;
    // rom_array[11941] = 32'h00009f49;
    // rom_array[11942] = 32'h00009f51;
    // rom_array[11943] = 32'hFFFFFFF0;
    // rom_array[11944] = 32'hFFFFFFF0;
    // rom_array[11945] = 32'h00009f59;
    // rom_array[11946] = 32'h00009f61;
    // rom_array[11947] = 32'h00009f69;
    // rom_array[11948] = 32'h00009f71;
    // rom_array[11949] = 32'hFFFFFFF0;
    // rom_array[11950] = 32'hFFFFFFF0;
    // rom_array[11951] = 32'hFFFFFFF0;
    // rom_array[11952] = 32'hFFFFFFF0;
    // rom_array[11953] = 32'h00009f79;
    // rom_array[11954] = 32'h00009f81;
    // rom_array[11955] = 32'h00009f89;
    // rom_array[11956] = 32'h00009f91;
    // rom_array[11957] = 32'hFFFFFFF0;
    // rom_array[11958] = 32'hFFFFFFF0;
    // rom_array[11959] = 32'hFFFFFFF0;
    // rom_array[11960] = 32'hFFFFFFF0;
    // rom_array[11961] = 32'h00009f99;
    // rom_array[11962] = 32'h00009fa1;
    // rom_array[11963] = 32'hFFFFFFF1;
    // rom_array[11964] = 32'hFFFFFFF1;
    // rom_array[11965] = 32'h00009fa9;
    // rom_array[11966] = 32'h00009fb1;
    // rom_array[11967] = 32'hFFFFFFF1;
    // rom_array[11968] = 32'hFFFFFFF1;
    // rom_array[11969] = 32'h00009fb9;
    // rom_array[11970] = 32'h00009fc1;
    // rom_array[11971] = 32'h00009fc9;
    // rom_array[11972] = 32'h00009fd1;
    // rom_array[11973] = 32'hFFFFFFF0;
    // rom_array[11974] = 32'hFFFFFFF0;
    // rom_array[11975] = 32'hFFFFFFF0;
    // rom_array[11976] = 32'hFFFFFFF0;
    // rom_array[11977] = 32'h00009fd9;
    // rom_array[11978] = 32'h00009fe1;
    // rom_array[11979] = 32'hFFFFFFF1;
    // rom_array[11980] = 32'hFFFFFFF1;
    // rom_array[11981] = 32'h00009fe9;
    // rom_array[11982] = 32'h00009ff1;
    // rom_array[11983] = 32'hFFFFFFF1;
    // rom_array[11984] = 32'hFFFFFFF1;
    // rom_array[11985] = 32'h00009ff9;
    // rom_array[11986] = 32'h0000a001;
    // rom_array[11987] = 32'hFFFFFFF1;
    // rom_array[11988] = 32'hFFFFFFF1;
    // rom_array[11989] = 32'h0000a009;
    // rom_array[11990] = 32'h0000a011;
    // rom_array[11991] = 32'hFFFFFFF1;
    // rom_array[11992] = 32'hFFFFFFF1;
    // rom_array[11993] = 32'h0000a019;
    // rom_array[11994] = 32'h0000a021;
    // rom_array[11995] = 32'hFFFFFFF1;
    // rom_array[11996] = 32'hFFFFFFF1;
    // rom_array[11997] = 32'h0000a029;
    // rom_array[11998] = 32'h0000a031;
    // rom_array[11999] = 32'h0000a039;
    // rom_array[12000] = 32'h0000a041;
    // rom_array[12001] = 32'h0000a049;
    // rom_array[12002] = 32'h0000a051;
    // rom_array[12003] = 32'hFFFFFFF0;
    // rom_array[12004] = 32'hFFFFFFF0;
    // rom_array[12005] = 32'h0000a059;
    // rom_array[12006] = 32'h0000a061;
    // rom_array[12007] = 32'hFFFFFFF0;
    // rom_array[12008] = 32'hFFFFFFF0;
    // rom_array[12009] = 32'h0000a069;
    // rom_array[12010] = 32'h0000a071;
    // rom_array[12011] = 32'hFFFFFFF0;
    // rom_array[12012] = 32'hFFFFFFF0;
    // rom_array[12013] = 32'h0000a079;
    // rom_array[12014] = 32'h0000a081;
    // rom_array[12015] = 32'hFFFFFFF0;
    // rom_array[12016] = 32'hFFFFFFF0;
    // rom_array[12017] = 32'h0000a089;
    // rom_array[12018] = 32'h0000a091;
    // rom_array[12019] = 32'hFFFFFFF0;
    // rom_array[12020] = 32'hFFFFFFF0;
    // rom_array[12021] = 32'h0000a099;
    // rom_array[12022] = 32'h0000a0a1;
    // rom_array[12023] = 32'hFFFFFFF0;
    // rom_array[12024] = 32'hFFFFFFF0;
    // rom_array[12025] = 32'hFFFFFFF1;
    // rom_array[12026] = 32'hFFFFFFF1;
    // rom_array[12027] = 32'hFFFFFFF1;
    // rom_array[12028] = 32'hFFFFFFF1;
    // rom_array[12029] = 32'h0000a0a9;
    // rom_array[12030] = 32'h0000a0b1;
    // rom_array[12031] = 32'h0000a0b9;
    // rom_array[12032] = 32'h0000a0c1;
    // rom_array[12033] = 32'h0000a0c9;
    // rom_array[12034] = 32'h0000a0d1;
    // rom_array[12035] = 32'hFFFFFFF0;
    // rom_array[12036] = 32'hFFFFFFF0;
    // rom_array[12037] = 32'h0000a0d9;
    // rom_array[12038] = 32'h0000a0e1;
    // rom_array[12039] = 32'hFFFFFFF0;
    // rom_array[12040] = 32'hFFFFFFF0;
    // rom_array[12041] = 32'h0000a0e9;
    // rom_array[12042] = 32'h0000a0f1;
    // rom_array[12043] = 32'h0000a0f9;
    // rom_array[12044] = 32'h0000a101;
    // rom_array[12045] = 32'hFFFFFFF1;
    // rom_array[12046] = 32'hFFFFFFF1;
    // rom_array[12047] = 32'hFFFFFFF1;
    // rom_array[12048] = 32'hFFFFFFF1;
    // rom_array[12049] = 32'h0000a109;
    // rom_array[12050] = 32'h0000a111;
    // rom_array[12051] = 32'h0000a119;
    // rom_array[12052] = 32'h0000a121;
    // rom_array[12053] = 32'hFFFFFFF1;
    // rom_array[12054] = 32'hFFFFFFF1;
    // rom_array[12055] = 32'hFFFFFFF1;
    // rom_array[12056] = 32'hFFFFFFF1;
    // rom_array[12057] = 32'h0000a129;
    // rom_array[12058] = 32'h0000a131;
    // rom_array[12059] = 32'h0000a139;
    // rom_array[12060] = 32'h0000a141;
    // rom_array[12061] = 32'hFFFFFFF1;
    // rom_array[12062] = 32'hFFFFFFF1;
    // rom_array[12063] = 32'hFFFFFFF1;
    // rom_array[12064] = 32'hFFFFFFF1;
    // rom_array[12065] = 32'h0000a149;
    // rom_array[12066] = 32'h0000a151;
    // rom_array[12067] = 32'h0000a159;
    // rom_array[12068] = 32'h0000a161;
    // rom_array[12069] = 32'hFFFFFFF1;
    // rom_array[12070] = 32'hFFFFFFF1;
    // rom_array[12071] = 32'hFFFFFFF1;
    // rom_array[12072] = 32'hFFFFFFF1;
    // rom_array[12073] = 32'h0000a169;
    // rom_array[12074] = 32'h0000a171;
    // rom_array[12075] = 32'h0000a179;
    // rom_array[12076] = 32'h0000a181;
    // rom_array[12077] = 32'hFFFFFFF1;
    // rom_array[12078] = 32'hFFFFFFF1;
    // rom_array[12079] = 32'hFFFFFFF1;
    // rom_array[12080] = 32'hFFFFFFF1;
    // rom_array[12081] = 32'h0000a189;
    // rom_array[12082] = 32'h0000a191;
    // rom_array[12083] = 32'hFFFFFFF0;
    // rom_array[12084] = 32'hFFFFFFF0;
    // rom_array[12085] = 32'h0000a199;
    // rom_array[12086] = 32'h0000a1a1;
    // rom_array[12087] = 32'hFFFFFFF0;
    // rom_array[12088] = 32'hFFFFFFF0;
    // rom_array[12089] = 32'h0000a1a9;
    // rom_array[12090] = 32'h0000a1b1;
    // rom_array[12091] = 32'hFFFFFFF0;
    // rom_array[12092] = 32'hFFFFFFF0;
    // rom_array[12093] = 32'h0000a1b9;
    // rom_array[12094] = 32'h0000a1c1;
    // rom_array[12095] = 32'hFFFFFFF0;
    // rom_array[12096] = 32'hFFFFFFF0;
    // rom_array[12097] = 32'h0000a1c9;
    // rom_array[12098] = 32'h0000a1d1;
    // rom_array[12099] = 32'hFFFFFFF0;
    // rom_array[12100] = 32'hFFFFFFF0;
    // rom_array[12101] = 32'h0000a1d9;
    // rom_array[12102] = 32'h0000a1e1;
    // rom_array[12103] = 32'hFFFFFFF0;
    // rom_array[12104] = 32'hFFFFFFF0;
    // rom_array[12105] = 32'h0000a1e9;
    // rom_array[12106] = 32'h0000a1f1;
    // rom_array[12107] = 32'hFFFFFFF0;
    // rom_array[12108] = 32'hFFFFFFF0;
    // rom_array[12109] = 32'h0000a1f9;
    // rom_array[12110] = 32'h0000a201;
    // rom_array[12111] = 32'hFFFFFFF0;
    // rom_array[12112] = 32'hFFFFFFF0;
    // rom_array[12113] = 32'h0000a209;
    // rom_array[12114] = 32'h0000a211;
    // rom_array[12115] = 32'h0000a219;
    // rom_array[12116] = 32'h0000a221;
    // rom_array[12117] = 32'hFFFFFFF1;
    // rom_array[12118] = 32'hFFFFFFF1;
    // rom_array[12119] = 32'hFFFFFFF1;
    // rom_array[12120] = 32'hFFFFFFF1;
    // rom_array[12121] = 32'h0000a229;
    // rom_array[12122] = 32'h0000a231;
    // rom_array[12123] = 32'h0000a239;
    // rom_array[12124] = 32'h0000a241;
    // rom_array[12125] = 32'hFFFFFFF1;
    // rom_array[12126] = 32'hFFFFFFF1;
    // rom_array[12127] = 32'hFFFFFFF1;
    // rom_array[12128] = 32'hFFFFFFF1;
    // rom_array[12129] = 32'h0000a249;
    // rom_array[12130] = 32'h0000a251;
    // rom_array[12131] = 32'h0000a259;
    // rom_array[12132] = 32'h0000a261;
    // rom_array[12133] = 32'hFFFFFFF1;
    // rom_array[12134] = 32'hFFFFFFF1;
    // rom_array[12135] = 32'hFFFFFFF1;
    // rom_array[12136] = 32'hFFFFFFF1;
    // rom_array[12137] = 32'h0000a269;
    // rom_array[12138] = 32'h0000a271;
    // rom_array[12139] = 32'h0000a279;
    // rom_array[12140] = 32'h0000a281;
    // rom_array[12141] = 32'h0000a289;
    // rom_array[12142] = 32'h0000a291;
    // rom_array[12143] = 32'hFFFFFFF1;
    // rom_array[12144] = 32'hFFFFFFF1;
    // rom_array[12145] = 32'h0000a299;
    // rom_array[12146] = 32'h0000a2a1;
    // rom_array[12147] = 32'hFFFFFFF1;
    // rom_array[12148] = 32'hFFFFFFF1;
    // rom_array[12149] = 32'h0000a2a9;
    // rom_array[12150] = 32'h0000a2b1;
    // rom_array[12151] = 32'hFFFFFFF1;
    // rom_array[12152] = 32'hFFFFFFF1;
    // rom_array[12153] = 32'h0000a2b9;
    // rom_array[12154] = 32'h0000a2c1;
    // rom_array[12155] = 32'h0000a2c9;
    // rom_array[12156] = 32'h0000a2d1;
    // rom_array[12157] = 32'hFFFFFFF0;
    // rom_array[12158] = 32'hFFFFFFF0;
    // rom_array[12159] = 32'hFFFFFFF0;
    // rom_array[12160] = 32'hFFFFFFF0;
    // rom_array[12161] = 32'h0000a2d9;
    // rom_array[12162] = 32'h0000a2e1;
    // rom_array[12163] = 32'h0000a2e9;
    // rom_array[12164] = 32'h0000a2f1;
    // rom_array[12165] = 32'hFFFFFFF0;
    // rom_array[12166] = 32'hFFFFFFF0;
    // rom_array[12167] = 32'hFFFFFFF0;
    // rom_array[12168] = 32'hFFFFFFF0;
    // rom_array[12169] = 32'h0000a2f9;
    // rom_array[12170] = 32'h0000a301;
    // rom_array[12171] = 32'h0000a309;
    // rom_array[12172] = 32'h0000a311;
    // rom_array[12173] = 32'hFFFFFFF0;
    // rom_array[12174] = 32'hFFFFFFF0;
    // rom_array[12175] = 32'hFFFFFFF0;
    // rom_array[12176] = 32'hFFFFFFF0;
    // rom_array[12177] = 32'h0000a319;
    // rom_array[12178] = 32'h0000a321;
    // rom_array[12179] = 32'h0000a329;
    // rom_array[12180] = 32'h0000a331;
    // rom_array[12181] = 32'hFFFFFFF0;
    // rom_array[12182] = 32'hFFFFFFF0;
    // rom_array[12183] = 32'hFFFFFFF0;
    // rom_array[12184] = 32'hFFFFFFF0;
    // rom_array[12185] = 32'h0000a339;
    // rom_array[12186] = 32'h0000a341;
    // rom_array[12187] = 32'h0000a349;
    // rom_array[12188] = 32'h0000a351;
    // rom_array[12189] = 32'hFFFFFFF1;
    // rom_array[12190] = 32'hFFFFFFF1;
    // rom_array[12191] = 32'hFFFFFFF1;
    // rom_array[12192] = 32'hFFFFFFF1;
    // rom_array[12193] = 32'h0000a359;
    // rom_array[12194] = 32'h0000a361;
    // rom_array[12195] = 32'hFFFFFFF0;
    // rom_array[12196] = 32'hFFFFFFF0;
    // rom_array[12197] = 32'h0000a369;
    // rom_array[12198] = 32'h0000a371;
    // rom_array[12199] = 32'hFFFFFFF0;
    // rom_array[12200] = 32'hFFFFFFF0;
    // rom_array[12201] = 32'h0000a379;
    // rom_array[12202] = 32'h0000a381;
    // rom_array[12203] = 32'hFFFFFFF0;
    // rom_array[12204] = 32'hFFFFFFF0;
    // rom_array[12205] = 32'h0000a389;
    // rom_array[12206] = 32'h0000a391;
    // rom_array[12207] = 32'hFFFFFFF0;
    // rom_array[12208] = 32'hFFFFFFF0;
    // rom_array[12209] = 32'h0000a399;
    // rom_array[12210] = 32'h0000a3a1;
    // rom_array[12211] = 32'h0000a3a9;
    // rom_array[12212] = 32'h0000a3b1;
    // rom_array[12213] = 32'hFFFFFFF0;
    // rom_array[12214] = 32'hFFFFFFF0;
    // rom_array[12215] = 32'hFFFFFFF0;
    // rom_array[12216] = 32'hFFFFFFF0;
    // rom_array[12217] = 32'h0000a3b9;
    // rom_array[12218] = 32'h0000a3c1;
    // rom_array[12219] = 32'hFFFFFFF0;
    // rom_array[12220] = 32'hFFFFFFF0;
    // rom_array[12221] = 32'h0000a3c9;
    // rom_array[12222] = 32'h0000a3d1;
    // rom_array[12223] = 32'hFFFFFFF0;
    // rom_array[12224] = 32'hFFFFFFF0;
    // rom_array[12225] = 32'h0000a3d9;
    // rom_array[12226] = 32'h0000a3e1;
    // rom_array[12227] = 32'hFFFFFFF0;
    // rom_array[12228] = 32'hFFFFFFF0;
    // rom_array[12229] = 32'h0000a3e9;
    // rom_array[12230] = 32'h0000a3f1;
    // rom_array[12231] = 32'hFFFFFFF0;
    // rom_array[12232] = 32'hFFFFFFF0;
    // rom_array[12233] = 32'h0000a3f9;
    // rom_array[12234] = 32'h0000a401;
    // rom_array[12235] = 32'h0000a409;
    // rom_array[12236] = 32'h0000a411;
    // rom_array[12237] = 32'hFFFFFFF0;
    // rom_array[12238] = 32'hFFFFFFF0;
    // rom_array[12239] = 32'hFFFFFFF0;
    // rom_array[12240] = 32'hFFFFFFF0;
    // rom_array[12241] = 32'h0000a419;
    // rom_array[12242] = 32'h0000a421;
    // rom_array[12243] = 32'h0000a429;
    // rom_array[12244] = 32'h0000a431;
    // rom_array[12245] = 32'hFFFFFFF0;
    // rom_array[12246] = 32'hFFFFFFF0;
    // rom_array[12247] = 32'hFFFFFFF0;
    // rom_array[12248] = 32'hFFFFFFF0;
    // rom_array[12249] = 32'h0000a439;
    // rom_array[12250] = 32'h0000a441;
    // rom_array[12251] = 32'h0000a449;
    // rom_array[12252] = 32'h0000a451;
    // rom_array[12253] = 32'hFFFFFFF0;
    // rom_array[12254] = 32'hFFFFFFF0;
    // rom_array[12255] = 32'hFFFFFFF0;
    // rom_array[12256] = 32'hFFFFFFF0;
    // rom_array[12257] = 32'h0000a459;
    // rom_array[12258] = 32'h0000a461;
    // rom_array[12259] = 32'h0000a469;
    // rom_array[12260] = 32'h0000a471;
    // rom_array[12261] = 32'hFFFFFFF0;
    // rom_array[12262] = 32'hFFFFFFF0;
    // rom_array[12263] = 32'hFFFFFFF0;
    // rom_array[12264] = 32'hFFFFFFF0;
    // rom_array[12265] = 32'h0000a479;
    // rom_array[12266] = 32'h0000a481;
    // rom_array[12267] = 32'hFFFFFFF0;
    // rom_array[12268] = 32'hFFFFFFF0;
    // rom_array[12269] = 32'h0000a489;
    // rom_array[12270] = 32'h0000a491;
    // rom_array[12271] = 32'hFFFFFFF0;
    // rom_array[12272] = 32'hFFFFFFF0;
    // rom_array[12273] = 32'h0000a499;
    // rom_array[12274] = 32'h0000a4a1;
    // rom_array[12275] = 32'hFFFFFFF0;
    // rom_array[12276] = 32'hFFFFFFF0;
    // rom_array[12277] = 32'h0000a4a9;
    // rom_array[12278] = 32'h0000a4b1;
    // rom_array[12279] = 32'hFFFFFFF0;
    // rom_array[12280] = 32'hFFFFFFF0;
    // rom_array[12281] = 32'h0000a4b9;
    // rom_array[12282] = 32'h0000a4c1;
    // rom_array[12283] = 32'h0000a4c9;
    // rom_array[12284] = 32'h0000a4d1;
    // rom_array[12285] = 32'hFFFFFFF0;
    // rom_array[12286] = 32'hFFFFFFF0;
    // rom_array[12287] = 32'hFFFFFFF0;
    // rom_array[12288] = 32'hFFFFFFF0;
    // rom_array[12289] = 32'h0000a4d9;
    // rom_array[12290] = 32'h0000a4e1;
    // rom_array[12291] = 32'hFFFFFFF0;
    // rom_array[12292] = 32'hFFFFFFF0;
    // rom_array[12293] = 32'hFFFFFFF0;
    // rom_array[12294] = 32'hFFFFFFF0;
    // rom_array[12295] = 32'hFFFFFFF0;
    // rom_array[12296] = 32'hFFFFFFF0;
    // rom_array[12297] = 32'h0000a4e9;
    // rom_array[12298] = 32'h0000a4f1;
    // rom_array[12299] = 32'h0000a4f9;
    // rom_array[12300] = 32'h0000a501;
    // rom_array[12301] = 32'hFFFFFFF1;
    // rom_array[12302] = 32'hFFFFFFF1;
    // rom_array[12303] = 32'hFFFFFFF1;
    // rom_array[12304] = 32'hFFFFFFF1;
    // rom_array[12305] = 32'h0000a509;
    // rom_array[12306] = 32'h0000a511;
    // rom_array[12307] = 32'h0000a519;
    // rom_array[12308] = 32'h0000a521;
    // rom_array[12309] = 32'hFFFFFFF1;
    // rom_array[12310] = 32'hFFFFFFF1;
    // rom_array[12311] = 32'hFFFFFFF1;
    // rom_array[12312] = 32'hFFFFFFF1;
    // rom_array[12313] = 32'h0000a529;
    // rom_array[12314] = 32'h0000a531;
    // rom_array[12315] = 32'h0000a539;
    // rom_array[12316] = 32'h0000a541;
    // rom_array[12317] = 32'hFFFFFFF1;
    // rom_array[12318] = 32'hFFFFFFF1;
    // rom_array[12319] = 32'hFFFFFFF1;
    // rom_array[12320] = 32'hFFFFFFF1;
    // rom_array[12321] = 32'h0000a549;
    // rom_array[12322] = 32'h0000a551;
    // rom_array[12323] = 32'h0000a559;
    // rom_array[12324] = 32'h0000a561;
    // rom_array[12325] = 32'hFFFFFFF1;
    // rom_array[12326] = 32'hFFFFFFF1;
    // rom_array[12327] = 32'hFFFFFFF1;
    // rom_array[12328] = 32'hFFFFFFF1;
    // rom_array[12329] = 32'h0000a569;
    // rom_array[12330] = 32'h0000a571;
    // rom_array[12331] = 32'h0000a579;
    // rom_array[12332] = 32'h0000a581;
    // rom_array[12333] = 32'hFFFFFFF1;
    // rom_array[12334] = 32'hFFFFFFF1;
    // rom_array[12335] = 32'hFFFFFFF1;
    // rom_array[12336] = 32'hFFFFFFF1;
    // rom_array[12337] = 32'h0000a589;
    // rom_array[12338] = 32'h0000a591;
    // rom_array[12339] = 32'hFFFFFFF0;
    // rom_array[12340] = 32'hFFFFFFF0;
    // rom_array[12341] = 32'h0000a599;
    // rom_array[12342] = 32'h0000a5a1;
    // rom_array[12343] = 32'hFFFFFFF0;
    // rom_array[12344] = 32'hFFFFFFF0;
    // rom_array[12345] = 32'h0000a5a9;
    // rom_array[12346] = 32'h0000a5b1;
    // rom_array[12347] = 32'hFFFFFFF0;
    // rom_array[12348] = 32'hFFFFFFF0;
    // rom_array[12349] = 32'h0000a5b9;
    // rom_array[12350] = 32'h0000a5c1;
    // rom_array[12351] = 32'hFFFFFFF0;
    // rom_array[12352] = 32'hFFFFFFF0;
    // rom_array[12353] = 32'h0000a5c9;
    // rom_array[12354] = 32'h0000a5d1;
    // rom_array[12355] = 32'h0000a5d9;
    // rom_array[12356] = 32'h0000a5e1;
    // rom_array[12357] = 32'hFFFFFFF0;
    // rom_array[12358] = 32'hFFFFFFF0;
    // rom_array[12359] = 32'hFFFFFFF0;
    // rom_array[12360] = 32'hFFFFFFF0;
    // rom_array[12361] = 32'h0000a5e9;
    // rom_array[12362] = 32'h0000a5f1;
    // rom_array[12363] = 32'h0000a5f9;
    // rom_array[12364] = 32'h0000a601;
    // rom_array[12365] = 32'hFFFFFFF0;
    // rom_array[12366] = 32'hFFFFFFF0;
    // rom_array[12367] = 32'hFFFFFFF0;
    // rom_array[12368] = 32'hFFFFFFF0;
    // rom_array[12369] = 32'h0000a609;
    // rom_array[12370] = 32'h0000a611;
    // rom_array[12371] = 32'h0000a619;
    // rom_array[12372] = 32'h0000a621;
    // rom_array[12373] = 32'hFFFFFFF0;
    // rom_array[12374] = 32'hFFFFFFF0;
    // rom_array[12375] = 32'hFFFFFFF0;
    // rom_array[12376] = 32'hFFFFFFF0;
    // rom_array[12377] = 32'h0000a629;
    // rom_array[12378] = 32'h0000a631;
    // rom_array[12379] = 32'h0000a639;
    // rom_array[12380] = 32'h0000a641;
    // rom_array[12381] = 32'hFFFFFFF0;
    // rom_array[12382] = 32'hFFFFFFF0;
    // rom_array[12383] = 32'hFFFFFFF0;
    // rom_array[12384] = 32'hFFFFFFF0;
    // rom_array[12385] = 32'h0000a649;
    // rom_array[12386] = 32'h0000a651;
    // rom_array[12387] = 32'h0000a659;
    // rom_array[12388] = 32'h0000a661;
    // rom_array[12389] = 32'hFFFFFFF0;
    // rom_array[12390] = 32'hFFFFFFF0;
    // rom_array[12391] = 32'hFFFFFFF0;
    // rom_array[12392] = 32'hFFFFFFF0;
    // rom_array[12393] = 32'h0000a669;
    // rom_array[12394] = 32'h0000a671;
    // rom_array[12395] = 32'hFFFFFFF0;
    // rom_array[12396] = 32'hFFFFFFF0;
    // rom_array[12397] = 32'hFFFFFFF0;
    // rom_array[12398] = 32'hFFFFFFF0;
    // rom_array[12399] = 32'hFFFFFFF0;
    // rom_array[12400] = 32'hFFFFFFF0;
    // rom_array[12401] = 32'h0000a679;
    // rom_array[12402] = 32'h0000a681;
    // rom_array[12403] = 32'h0000a689;
    // rom_array[12404] = 32'h0000a691;
    // rom_array[12405] = 32'hFFFFFFF0;
    // rom_array[12406] = 32'hFFFFFFF0;
    // rom_array[12407] = 32'hFFFFFFF0;
    // rom_array[12408] = 32'hFFFFFFF0;
    // rom_array[12409] = 32'h0000a699;
    // rom_array[12410] = 32'h0000a6a1;
    // rom_array[12411] = 32'h0000a6a9;
    // rom_array[12412] = 32'h0000a6b1;
    // rom_array[12413] = 32'hFFFFFFF0;
    // rom_array[12414] = 32'hFFFFFFF0;
    // rom_array[12415] = 32'hFFFFFFF0;
    // rom_array[12416] = 32'hFFFFFFF0;
    // rom_array[12417] = 32'h0000a6b9;
    // rom_array[12418] = 32'h0000a6c1;
    // rom_array[12419] = 32'h0000a6c9;
    // rom_array[12420] = 32'h0000a6d1;
    // rom_array[12421] = 32'hFFFFFFF0;
    // rom_array[12422] = 32'hFFFFFFF0;
    // rom_array[12423] = 32'hFFFFFFF0;
    // rom_array[12424] = 32'hFFFFFFF0;
    // rom_array[12425] = 32'h0000a6d9;
    // rom_array[12426] = 32'h0000a6e1;
    // rom_array[12427] = 32'hFFFFFFF0;
    // rom_array[12428] = 32'hFFFFFFF0;
    // rom_array[12429] = 32'hFFFFFFF0;
    // rom_array[12430] = 32'hFFFFFFF0;
    // rom_array[12431] = 32'hFFFFFFF0;
    // rom_array[12432] = 32'hFFFFFFF0;
    // rom_array[12433] = 32'h0000a6e9;
    // rom_array[12434] = 32'h0000a6f1;
    // rom_array[12435] = 32'h0000a6f9;
    // rom_array[12436] = 32'h0000a701;
    // rom_array[12437] = 32'hFFFFFFF1;
    // rom_array[12438] = 32'hFFFFFFF1;
    // rom_array[12439] = 32'hFFFFFFF1;
    // rom_array[12440] = 32'hFFFFFFF1;
    // rom_array[12441] = 32'h0000a709;
    // rom_array[12442] = 32'h0000a711;
    // rom_array[12443] = 32'h0000a719;
    // rom_array[12444] = 32'h0000a721;
    // rom_array[12445] = 32'hFFFFFFF1;
    // rom_array[12446] = 32'hFFFFFFF1;
    // rom_array[12447] = 32'hFFFFFFF1;
    // rom_array[12448] = 32'hFFFFFFF1;
    // rom_array[12449] = 32'h0000a729;
    // rom_array[12450] = 32'h0000a731;
    // rom_array[12451] = 32'h0000a739;
    // rom_array[12452] = 32'h0000a741;
    // rom_array[12453] = 32'hFFFFFFF1;
    // rom_array[12454] = 32'hFFFFFFF1;
    // rom_array[12455] = 32'hFFFFFFF1;
    // rom_array[12456] = 32'hFFFFFFF1;
    // rom_array[12457] = 32'h0000a749;
    // rom_array[12458] = 32'h0000a751;
    // rom_array[12459] = 32'h0000a759;
    // rom_array[12460] = 32'h0000a761;
    // rom_array[12461] = 32'hFFFFFFF1;
    // rom_array[12462] = 32'hFFFFFFF1;
    // rom_array[12463] = 32'hFFFFFFF1;
    // rom_array[12464] = 32'hFFFFFFF1;
    // rom_array[12465] = 32'h0000a769;
    // rom_array[12466] = 32'h0000a771;
    // rom_array[12467] = 32'h0000a779;
    // rom_array[12468] = 32'h0000a781;
    // rom_array[12469] = 32'h0000a789;
    // rom_array[12470] = 32'h0000a791;
    // rom_array[12471] = 32'hFFFFFFF0;
    // rom_array[12472] = 32'hFFFFFFF0;
    // rom_array[12473] = 32'h0000a799;
    // rom_array[12474] = 32'h0000a7a1;
    // rom_array[12475] = 32'h0000a7a9;
    // rom_array[12476] = 32'h0000a7b1;
    // rom_array[12477] = 32'hFFFFFFF0;
    // rom_array[12478] = 32'hFFFFFFF0;
    // rom_array[12479] = 32'hFFFFFFF0;
    // rom_array[12480] = 32'hFFFFFFF0;
    // rom_array[12481] = 32'h0000a7b9;
    // rom_array[12482] = 32'h0000a7c1;
    // rom_array[12483] = 32'h0000a7c9;
    // rom_array[12484] = 32'h0000a7d1;
    // rom_array[12485] = 32'hFFFFFFF0;
    // rom_array[12486] = 32'hFFFFFFF0;
    // rom_array[12487] = 32'hFFFFFFF0;
    // rom_array[12488] = 32'hFFFFFFF0;
    // rom_array[12489] = 32'h0000a7d9;
    // rom_array[12490] = 32'h0000a7e1;
    // rom_array[12491] = 32'h0000a7e9;
    // rom_array[12492] = 32'h0000a7f1;
    // rom_array[12493] = 32'h0000a7f9;
    // rom_array[12494] = 32'h0000a801;
    // rom_array[12495] = 32'hFFFFFFF1;
    // rom_array[12496] = 32'hFFFFFFF1;
    // rom_array[12497] = 32'h0000a809;
    // rom_array[12498] = 32'h0000a811;
    // rom_array[12499] = 32'h0000a819;
    // rom_array[12500] = 32'h0000a821;
    // rom_array[12501] = 32'hFFFFFFF1;
    // rom_array[12502] = 32'hFFFFFFF1;
    // rom_array[12503] = 32'hFFFFFFF1;
    // rom_array[12504] = 32'hFFFFFFF1;
    // rom_array[12505] = 32'h0000a829;
    // rom_array[12506] = 32'h0000a831;
    // rom_array[12507] = 32'hFFFFFFF0;
    // rom_array[12508] = 32'hFFFFFFF0;
    // rom_array[12509] = 32'h0000a839;
    // rom_array[12510] = 32'h0000a841;
    // rom_array[12511] = 32'hFFFFFFF0;
    // rom_array[12512] = 32'hFFFFFFF0;
    // rom_array[12513] = 32'h0000a849;
    // rom_array[12514] = 32'h0000a851;
    // rom_array[12515] = 32'hFFFFFFF0;
    // rom_array[12516] = 32'hFFFFFFF0;
    // rom_array[12517] = 32'h0000a859;
    // rom_array[12518] = 32'h0000a861;
    // rom_array[12519] = 32'hFFFFFFF0;
    // rom_array[12520] = 32'hFFFFFFF0;
    // rom_array[12521] = 32'h0000a869;
    // rom_array[12522] = 32'h0000a871;
    // rom_array[12523] = 32'h0000a879;
    // rom_array[12524] = 32'h0000a881;
    // rom_array[12525] = 32'hFFFFFFF1;
    // rom_array[12526] = 32'hFFFFFFF1;
    // rom_array[12527] = 32'hFFFFFFF1;
    // rom_array[12528] = 32'hFFFFFFF1;
    // rom_array[12529] = 32'h0000a889;
    // rom_array[12530] = 32'h0000a891;
    // rom_array[12531] = 32'hFFFFFFF0;
    // rom_array[12532] = 32'hFFFFFFF0;
    // rom_array[12533] = 32'h0000a899;
    // rom_array[12534] = 32'h0000a8a1;
    // rom_array[12535] = 32'hFFFFFFF0;
    // rom_array[12536] = 32'hFFFFFFF0;
    // rom_array[12537] = 32'h0000a8a9;
    // rom_array[12538] = 32'h0000a8b1;
    // rom_array[12539] = 32'hFFFFFFF0;
    // rom_array[12540] = 32'hFFFFFFF0;
    // rom_array[12541] = 32'h0000a8b9;
    // rom_array[12542] = 32'h0000a8c1;
    // rom_array[12543] = 32'hFFFFFFF0;
    // rom_array[12544] = 32'hFFFFFFF0;
    // rom_array[12545] = 32'h0000a8c9;
    // rom_array[12546] = 32'h0000a8d1;
    // rom_array[12547] = 32'hFFFFFFF0;
    // rom_array[12548] = 32'hFFFFFFF0;
    // rom_array[12549] = 32'h0000a8d9;
    // rom_array[12550] = 32'h0000a8e1;
    // rom_array[12551] = 32'hFFFFFFF0;
    // rom_array[12552] = 32'hFFFFFFF0;
    // rom_array[12553] = 32'h0000a8e9;
    // rom_array[12554] = 32'h0000a8f1;
    // rom_array[12555] = 32'hFFFFFFF1;
    // rom_array[12556] = 32'hFFFFFFF1;
    // rom_array[12557] = 32'h0000a8f9;
    // rom_array[12558] = 32'h0000a901;
    // rom_array[12559] = 32'hFFFFFFF1;
    // rom_array[12560] = 32'hFFFFFFF1;
    // rom_array[12561] = 32'h0000a909;
    // rom_array[12562] = 32'h0000a911;
    // rom_array[12563] = 32'hFFFFFFF1;
    // rom_array[12564] = 32'hFFFFFFF1;
    // rom_array[12565] = 32'h0000a919;
    // rom_array[12566] = 32'h0000a921;
    // rom_array[12567] = 32'hFFFFFFF1;
    // rom_array[12568] = 32'hFFFFFFF1;
    // rom_array[12569] = 32'h0000a929;
    // rom_array[12570] = 32'h0000a931;
    // rom_array[12571] = 32'hFFFFFFF0;
    // rom_array[12572] = 32'hFFFFFFF0;
    // rom_array[12573] = 32'h0000a939;
    // rom_array[12574] = 32'h0000a941;
    // rom_array[12575] = 32'h0000a949;
    // rom_array[12576] = 32'h0000a951;
    // rom_array[12577] = 32'hFFFFFFF0;
    // rom_array[12578] = 32'hFFFFFFF0;
    // rom_array[12579] = 32'hFFFFFFF0;
    // rom_array[12580] = 32'hFFFFFFF0;
    // rom_array[12581] = 32'h0000a959;
    // rom_array[12582] = 32'h0000a961;
    // rom_array[12583] = 32'h0000a969;
    // rom_array[12584] = 32'h0000a971;
    // rom_array[12585] = 32'h0000a979;
    // rom_array[12586] = 32'h0000a981;
    // rom_array[12587] = 32'hFFFFFFF0;
    // rom_array[12588] = 32'hFFFFFFF0;
    // rom_array[12589] = 32'hFFFFFFF0;
    // rom_array[12590] = 32'hFFFFFFF0;
    // rom_array[12591] = 32'hFFFFFFF0;
    // rom_array[12592] = 32'hFFFFFFF0;
    // rom_array[12593] = 32'hFFFFFFF0;
    // rom_array[12594] = 32'hFFFFFFF0;
    // rom_array[12595] = 32'hFFFFFFF0;
    // rom_array[12596] = 32'hFFFFFFF0;
    // rom_array[12597] = 32'h0000a989;
    // rom_array[12598] = 32'h0000a991;
    // rom_array[12599] = 32'h0000a999;
    // rom_array[12600] = 32'h0000a9a1;
    // rom_array[12601] = 32'h0000a9a9;
    // rom_array[12602] = 32'h0000a9b1;
    // rom_array[12603] = 32'hFFFFFFF1;
    // rom_array[12604] = 32'hFFFFFFF1;
    // rom_array[12605] = 32'h0000a9b9;
    // rom_array[12606] = 32'h0000a9c1;
    // rom_array[12607] = 32'h0000a9c9;
    // rom_array[12608] = 32'h0000a9d1;
    // rom_array[12609] = 32'h0000a9d9;
    // rom_array[12610] = 32'h0000a9e1;
    // rom_array[12611] = 32'h0000a9e9;
    // rom_array[12612] = 32'h0000a9f1;
    // rom_array[12613] = 32'hFFFFFFF1;
    // rom_array[12614] = 32'hFFFFFFF1;
    // rom_array[12615] = 32'h0000a9f9;
    // rom_array[12616] = 32'h0000aa01;
    // rom_array[12617] = 32'h0000aa09;
    // rom_array[12618] = 32'h0000aa11;
    // rom_array[12619] = 32'hFFFFFFF0;
    // rom_array[12620] = 32'hFFFFFFF0;
    // rom_array[12621] = 32'h0000aa19;
    // rom_array[12622] = 32'h0000aa21;
    // rom_array[12623] = 32'hFFFFFFF0;
    // rom_array[12624] = 32'hFFFFFFF0;
    // rom_array[12625] = 32'h0000aa29;
    // rom_array[12626] = 32'h0000aa31;
    // rom_array[12627] = 32'hFFFFFFF0;
    // rom_array[12628] = 32'hFFFFFFF0;
    // rom_array[12629] = 32'h0000aa39;
    // rom_array[12630] = 32'h0000aa41;
    // rom_array[12631] = 32'hFFFFFFF0;
    // rom_array[12632] = 32'hFFFFFFF0;
    // rom_array[12633] = 32'h0000aa49;
    // rom_array[12634] = 32'h0000aa51;
    // rom_array[12635] = 32'hFFFFFFF0;
    // rom_array[12636] = 32'hFFFFFFF0;
    // rom_array[12637] = 32'h0000aa59;
    // rom_array[12638] = 32'h0000aa61;
    // rom_array[12639] = 32'hFFFFFFF0;
    // rom_array[12640] = 32'hFFFFFFF0;
    // rom_array[12641] = 32'h0000aa69;
    // rom_array[12642] = 32'h0000aa71;
    // rom_array[12643] = 32'h0000aa79;
    // rom_array[12644] = 32'h0000aa81;
    // rom_array[12645] = 32'hFFFFFFF0;
    // rom_array[12646] = 32'hFFFFFFF0;
    // rom_array[12647] = 32'hFFFFFFF0;
    // rom_array[12648] = 32'hFFFFFFF0;
    // rom_array[12649] = 32'h0000aa89;
    // rom_array[12650] = 32'h0000aa91;
    // rom_array[12651] = 32'hFFFFFFF0;
    // rom_array[12652] = 32'hFFFFFFF0;
    // rom_array[12653] = 32'hFFFFFFF0;
    // rom_array[12654] = 32'hFFFFFFF0;
    // rom_array[12655] = 32'hFFFFFFF0;
    // rom_array[12656] = 32'hFFFFFFF0;
    // rom_array[12657] = 32'hFFFFFFF1;
    // rom_array[12658] = 32'hFFFFFFF1;
    // rom_array[12659] = 32'hFFFFFFF1;
    // rom_array[12660] = 32'hFFFFFFF1;
    // rom_array[12661] = 32'h0000aa99;
    // rom_array[12662] = 32'h0000aaa1;
    // rom_array[12663] = 32'h0000aaa9;
    // rom_array[12664] = 32'h0000aab1;
    // rom_array[12665] = 32'hFFFFFFF1;
    // rom_array[12666] = 32'hFFFFFFF1;
    // rom_array[12667] = 32'hFFFFFFF1;
    // rom_array[12668] = 32'hFFFFFFF1;
    // rom_array[12669] = 32'h0000aab9;
    // rom_array[12670] = 32'h0000aac1;
    // rom_array[12671] = 32'h0000aac9;
    // rom_array[12672] = 32'h0000aad1;
    // rom_array[12673] = 32'hFFFFFFF1;
    // rom_array[12674] = 32'hFFFFFFF1;
    // rom_array[12675] = 32'hFFFFFFF1;
    // rom_array[12676] = 32'hFFFFFFF1;
    // rom_array[12677] = 32'h0000aad9;
    // rom_array[12678] = 32'h0000aae1;
    // rom_array[12679] = 32'h0000aae9;
    // rom_array[12680] = 32'h0000aaf1;
    // rom_array[12681] = 32'hFFFFFFF1;
    // rom_array[12682] = 32'hFFFFFFF1;
    // rom_array[12683] = 32'h0000aaf9;
    // rom_array[12684] = 32'h0000ab01;
    // rom_array[12685] = 32'h0000ab09;
    // rom_array[12686] = 32'h0000ab11;
    // rom_array[12687] = 32'h0000ab19;
    // rom_array[12688] = 32'h0000ab21;
    // rom_array[12689] = 32'hFFFFFFF0;
    // rom_array[12690] = 32'hFFFFFFF0;
    // rom_array[12691] = 32'hFFFFFFF0;
    // rom_array[12692] = 32'hFFFFFFF0;
    // rom_array[12693] = 32'h0000ab29;
    // rom_array[12694] = 32'h0000ab31;
    // rom_array[12695] = 32'h0000ab39;
    // rom_array[12696] = 32'h0000ab41;
    // rom_array[12697] = 32'h0000ab49;
    // rom_array[12698] = 32'h0000ab51;
    // rom_array[12699] = 32'hFFFFFFF1;
    // rom_array[12700] = 32'hFFFFFFF1;
    // rom_array[12701] = 32'h0000ab59;
    // rom_array[12702] = 32'h0000ab61;
    // rom_array[12703] = 32'hFFFFFFF1;
    // rom_array[12704] = 32'hFFFFFFF1;
    // rom_array[12705] = 32'h0000ab69;
    // rom_array[12706] = 32'h0000ab71;
    // rom_array[12707] = 32'h0000ab79;
    // rom_array[12708] = 32'h0000ab81;
    // rom_array[12709] = 32'hFFFFFFF1;
    // rom_array[12710] = 32'hFFFFFFF1;
    // rom_array[12711] = 32'hFFFFFFF1;
    // rom_array[12712] = 32'hFFFFFFF1;
    // rom_array[12713] = 32'h0000ab89;
    // rom_array[12714] = 32'h0000ab91;
    // rom_array[12715] = 32'h0000ab99;
    // rom_array[12716] = 32'h0000aba1;
    // rom_array[12717] = 32'hFFFFFFF1;
    // rom_array[12718] = 32'hFFFFFFF1;
    // rom_array[12719] = 32'hFFFFFFF1;
    // rom_array[12720] = 32'hFFFFFFF1;
    // rom_array[12721] = 32'h0000aba9;
    // rom_array[12722] = 32'h0000abb1;
    // rom_array[12723] = 32'hFFFFFFF1;
    // rom_array[12724] = 32'hFFFFFFF1;
    // rom_array[12725] = 32'h0000abb9;
    // rom_array[12726] = 32'h0000abc1;
    // rom_array[12727] = 32'hFFFFFFF1;
    // rom_array[12728] = 32'hFFFFFFF1;
    // rom_array[12729] = 32'h0000abc9;
    // rom_array[12730] = 32'h0000abd1;
    // rom_array[12731] = 32'h0000abd9;
    // rom_array[12732] = 32'h0000abe1;
    // rom_array[12733] = 32'hFFFFFFF1;
    // rom_array[12734] = 32'hFFFFFFF1;
    // rom_array[12735] = 32'hFFFFFFF1;
    // rom_array[12736] = 32'hFFFFFFF1;
    // rom_array[12737] = 32'h0000abe9;
    // rom_array[12738] = 32'h0000abf1;
    // rom_array[12739] = 32'hFFFFFFF1;
    // rom_array[12740] = 32'hFFFFFFF1;
    // rom_array[12741] = 32'h0000abf9;
    // rom_array[12742] = 32'h0000ac01;
    // rom_array[12743] = 32'hFFFFFFF1;
    // rom_array[12744] = 32'hFFFFFFF1;
    // rom_array[12745] = 32'hFFFFFFF0;
    // rom_array[12746] = 32'hFFFFFFF0;
    // rom_array[12747] = 32'hFFFFFFF0;
    // rom_array[12748] = 32'hFFFFFFF0;
    // rom_array[12749] = 32'h0000ac09;
    // rom_array[12750] = 32'h0000ac11;
    // rom_array[12751] = 32'h0000ac19;
    // rom_array[12752] = 32'h0000ac21;
    // rom_array[12753] = 32'hFFFFFFF0;
    // rom_array[12754] = 32'hFFFFFFF0;
    // rom_array[12755] = 32'hFFFFFFF0;
    // rom_array[12756] = 32'hFFFFFFF0;
    // rom_array[12757] = 32'h0000ac29;
    // rom_array[12758] = 32'h0000ac31;
    // rom_array[12759] = 32'hFFFFFFF0;
    // rom_array[12760] = 32'hFFFFFFF0;
    // rom_array[12761] = 32'h0000ac39;
    // rom_array[12762] = 32'h0000ac41;
    // rom_array[12763] = 32'hFFFFFFF0;
    // rom_array[12764] = 32'hFFFFFFF0;
    // rom_array[12765] = 32'h0000ac49;
    // rom_array[12766] = 32'h0000ac51;
    // rom_array[12767] = 32'hFFFFFFF0;
    // rom_array[12768] = 32'hFFFFFFF0;
    // rom_array[12769] = 32'h0000ac59;
    // rom_array[12770] = 32'h0000ac61;
    // rom_array[12771] = 32'hFFFFFFF0;
    // rom_array[12772] = 32'hFFFFFFF0;
    // rom_array[12773] = 32'h0000ac69;
    // rom_array[12774] = 32'h0000ac71;
    // rom_array[12775] = 32'hFFFFFFF0;
    // rom_array[12776] = 32'hFFFFFFF0;
    // rom_array[12777] = 32'h0000ac79;
    // rom_array[12778] = 32'h0000ac81;
    // rom_array[12779] = 32'hFFFFFFF0;
    // rom_array[12780] = 32'hFFFFFFF0;
    // rom_array[12781] = 32'h0000ac89;
    // rom_array[12782] = 32'h0000ac91;
    // rom_array[12783] = 32'hFFFFFFF0;
    // rom_array[12784] = 32'hFFFFFFF0;
    // rom_array[12785] = 32'h0000ac99;
    // rom_array[12786] = 32'h0000aca1;
    // rom_array[12787] = 32'h0000aca9;
    // rom_array[12788] = 32'h0000acb1;
    // rom_array[12789] = 32'hFFFFFFF0;
    // rom_array[12790] = 32'hFFFFFFF0;
    // rom_array[12791] = 32'hFFFFFFF0;
    // rom_array[12792] = 32'hFFFFFFF0;
    // rom_array[12793] = 32'h0000acb9;
    // rom_array[12794] = 32'h0000acc1;
    // rom_array[12795] = 32'h0000acc9;
    // rom_array[12796] = 32'h0000acd1;
    // rom_array[12797] = 32'hFFFFFFF0;
    // rom_array[12798] = 32'hFFFFFFF0;
    // rom_array[12799] = 32'hFFFFFFF0;
    // rom_array[12800] = 32'hFFFFFFF0;
    // rom_array[12801] = 32'h0000acd9;
    // rom_array[12802] = 32'h0000ace1;
    // rom_array[12803] = 32'hFFFFFFF1;
    // rom_array[12804] = 32'hFFFFFFF1;
    // rom_array[12805] = 32'h0000ace9;
    // rom_array[12806] = 32'h0000acf1;
    // rom_array[12807] = 32'hFFFFFFF1;
    // rom_array[12808] = 32'hFFFFFFF1;
    // rom_array[12809] = 32'h0000acf9;
    // rom_array[12810] = 32'h0000ad01;
    // rom_array[12811] = 32'h0000ad09;
    // rom_array[12812] = 32'h0000ad11;
    // rom_array[12813] = 32'hFFFFFFF0;
    // rom_array[12814] = 32'hFFFFFFF0;
    // rom_array[12815] = 32'hFFFFFFF0;
    // rom_array[12816] = 32'hFFFFFFF0;
    // rom_array[12817] = 32'h0000ad19;
    // rom_array[12818] = 32'h0000ad21;
    // rom_array[12819] = 32'hFFFFFFF1;
    // rom_array[12820] = 32'hFFFFFFF1;
    // rom_array[12821] = 32'h0000ad29;
    // rom_array[12822] = 32'h0000ad31;
    // rom_array[12823] = 32'hFFFFFFF1;
    // rom_array[12824] = 32'hFFFFFFF1;
    // rom_array[12825] = 32'h0000ad39;
    // rom_array[12826] = 32'h0000ad41;
    // rom_array[12827] = 32'hFFFFFFF1;
    // rom_array[12828] = 32'hFFFFFFF1;
    // rom_array[12829] = 32'h0000ad49;
    // rom_array[12830] = 32'h0000ad51;
    // rom_array[12831] = 32'hFFFFFFF1;
    // rom_array[12832] = 32'hFFFFFFF1;
    // rom_array[12833] = 32'h0000ad59;
    // rom_array[12834] = 32'h0000ad61;
    // rom_array[12835] = 32'hFFFFFFF1;
    // rom_array[12836] = 32'hFFFFFFF1;
    // rom_array[12837] = 32'h0000ad69;
    // rom_array[12838] = 32'h0000ad71;
    // rom_array[12839] = 32'h0000ad79;
    // rom_array[12840] = 32'h0000ad81;
    // rom_array[12841] = 32'h0000ad89;
    // rom_array[12842] = 32'h0000ad91;
    // rom_array[12843] = 32'hFFFFFFF0;
    // rom_array[12844] = 32'hFFFFFFF0;
    // rom_array[12845] = 32'h0000ad99;
    // rom_array[12846] = 32'h0000ada1;
    // rom_array[12847] = 32'hFFFFFFF0;
    // rom_array[12848] = 32'hFFFFFFF0;
    // rom_array[12849] = 32'h0000ada9;
    // rom_array[12850] = 32'h0000adb1;
    // rom_array[12851] = 32'hFFFFFFF0;
    // rom_array[12852] = 32'hFFFFFFF0;
    // rom_array[12853] = 32'h0000adb9;
    // rom_array[12854] = 32'h0000adc1;
    // rom_array[12855] = 32'hFFFFFFF0;
    // rom_array[12856] = 32'hFFFFFFF0;
    // rom_array[12857] = 32'h0000adc9;
    // rom_array[12858] = 32'h0000add1;
    // rom_array[12859] = 32'hFFFFFFF0;
    // rom_array[12860] = 32'hFFFFFFF0;
    // rom_array[12861] = 32'h0000add9;
    // rom_array[12862] = 32'h0000ade1;
    // rom_array[12863] = 32'hFFFFFFF0;
    // rom_array[12864] = 32'hFFFFFFF0;
    // rom_array[12865] = 32'hFFFFFFF1;
    // rom_array[12866] = 32'hFFFFFFF1;
    // rom_array[12867] = 32'hFFFFFFF1;
    // rom_array[12868] = 32'hFFFFFFF1;
    // rom_array[12869] = 32'h0000ade9;
    // rom_array[12870] = 32'h0000adf1;
    // rom_array[12871] = 32'h0000adf9;
    // rom_array[12872] = 32'h0000ae01;
    // rom_array[12873] = 32'h0000ae09;
    // rom_array[12874] = 32'h0000ae11;
    // rom_array[12875] = 32'hFFFFFFF0;
    // rom_array[12876] = 32'hFFFFFFF0;
    // rom_array[12877] = 32'h0000ae19;
    // rom_array[12878] = 32'h0000ae21;
    // rom_array[12879] = 32'hFFFFFFF0;
    // rom_array[12880] = 32'hFFFFFFF0;
    // rom_array[12881] = 32'h0000ae29;
    // rom_array[12882] = 32'h0000ae31;
    // rom_array[12883] = 32'h0000ae39;
    // rom_array[12884] = 32'h0000ae41;
    // rom_array[12885] = 32'hFFFFFFF1;
    // rom_array[12886] = 32'hFFFFFFF1;
    // rom_array[12887] = 32'hFFFFFFF1;
    // rom_array[12888] = 32'hFFFFFFF1;
    // rom_array[12889] = 32'h0000ae49;
    // rom_array[12890] = 32'h0000ae51;
    // rom_array[12891] = 32'h0000ae59;
    // rom_array[12892] = 32'h0000ae61;
    // rom_array[12893] = 32'hFFFFFFF1;
    // rom_array[12894] = 32'hFFFFFFF1;
    // rom_array[12895] = 32'hFFFFFFF1;
    // rom_array[12896] = 32'hFFFFFFF1;
    // rom_array[12897] = 32'h0000ae69;
    // rom_array[12898] = 32'h0000ae71;
    // rom_array[12899] = 32'h0000ae79;
    // rom_array[12900] = 32'h0000ae81;
    // rom_array[12901] = 32'hFFFFFFF1;
    // rom_array[12902] = 32'hFFFFFFF1;
    // rom_array[12903] = 32'hFFFFFFF1;
    // rom_array[12904] = 32'hFFFFFFF1;
    // rom_array[12905] = 32'h0000ae89;
    // rom_array[12906] = 32'h0000ae91;
    // rom_array[12907] = 32'h0000ae99;
    // rom_array[12908] = 32'h0000aea1;
    // rom_array[12909] = 32'hFFFFFFF1;
    // rom_array[12910] = 32'hFFFFFFF1;
    // rom_array[12911] = 32'hFFFFFFF1;
    // rom_array[12912] = 32'hFFFFFFF1;
    // rom_array[12913] = 32'h0000aea9;
    // rom_array[12914] = 32'h0000aeb1;
    // rom_array[12915] = 32'h0000aeb9;
    // rom_array[12916] = 32'h0000aec1;
    // rom_array[12917] = 32'hFFFFFFF1;
    // rom_array[12918] = 32'hFFFFFFF1;
    // rom_array[12919] = 32'hFFFFFFF1;
    // rom_array[12920] = 32'hFFFFFFF1;
    // rom_array[12921] = 32'h0000aec9;
    // rom_array[12922] = 32'h0000aed1;
    // rom_array[12923] = 32'hFFFFFFF0;
    // rom_array[12924] = 32'hFFFFFFF0;
    // rom_array[12925] = 32'h0000aed9;
    // rom_array[12926] = 32'h0000aee1;
    // rom_array[12927] = 32'hFFFFFFF0;
    // rom_array[12928] = 32'hFFFFFFF0;
    // rom_array[12929] = 32'h0000aee9;
    // rom_array[12930] = 32'h0000aef1;
    // rom_array[12931] = 32'hFFFFFFF0;
    // rom_array[12932] = 32'hFFFFFFF0;
    // rom_array[12933] = 32'h0000aef9;
    // rom_array[12934] = 32'h0000af01;
    // rom_array[12935] = 32'hFFFFFFF0;
    // rom_array[12936] = 32'hFFFFFFF0;
    // rom_array[12937] = 32'h0000af09;
    // rom_array[12938] = 32'h0000af11;
    // rom_array[12939] = 32'hFFFFFFF0;
    // rom_array[12940] = 32'hFFFFFFF0;
    // rom_array[12941] = 32'h0000af19;
    // rom_array[12942] = 32'h0000af21;
    // rom_array[12943] = 32'hFFFFFFF0;
    // rom_array[12944] = 32'hFFFFFFF0;
    // rom_array[12945] = 32'h0000af29;
    // rom_array[12946] = 32'h0000af31;
    // rom_array[12947] = 32'hFFFFFFF0;
    // rom_array[12948] = 32'hFFFFFFF0;
    // rom_array[12949] = 32'h0000af39;
    // rom_array[12950] = 32'h0000af41;
    // rom_array[12951] = 32'hFFFFFFF0;
    // rom_array[12952] = 32'hFFFFFFF0;
    // rom_array[12953] = 32'h0000af49;
    // rom_array[12954] = 32'h0000af51;
    // rom_array[12955] = 32'h0000af59;
    // rom_array[12956] = 32'h0000af61;
    // rom_array[12957] = 32'hFFFFFFF1;
    // rom_array[12958] = 32'hFFFFFFF1;
    // rom_array[12959] = 32'hFFFFFFF1;
    // rom_array[12960] = 32'hFFFFFFF1;
    // rom_array[12961] = 32'h0000af69;
    // rom_array[12962] = 32'h0000af71;
    // rom_array[12963] = 32'h0000af79;
    // rom_array[12964] = 32'h0000af81;
    // rom_array[12965] = 32'hFFFFFFF1;
    // rom_array[12966] = 32'hFFFFFFF1;
    // rom_array[12967] = 32'hFFFFFFF1;
    // rom_array[12968] = 32'hFFFFFFF1;
    // rom_array[12969] = 32'h0000af89;
    // rom_array[12970] = 32'h0000af91;
    // rom_array[12971] = 32'h0000af99;
    // rom_array[12972] = 32'h0000afa1;
    // rom_array[12973] = 32'hFFFFFFF1;
    // rom_array[12974] = 32'hFFFFFFF1;
    // rom_array[12975] = 32'hFFFFFFF1;
    // rom_array[12976] = 32'hFFFFFFF1;
    // rom_array[12977] = 32'h0000afa9;
    // rom_array[12978] = 32'h0000afb1;
    // rom_array[12979] = 32'h0000afb9;
    // rom_array[12980] = 32'h0000afc1;
    // rom_array[12981] = 32'h0000afc9;
    // rom_array[12982] = 32'h0000afd1;
    // rom_array[12983] = 32'hFFFFFFF1;
    // rom_array[12984] = 32'hFFFFFFF1;
    // rom_array[12985] = 32'h0000afd9;
    // rom_array[12986] = 32'h0000afe1;
    // rom_array[12987] = 32'hFFFFFFF1;
    // rom_array[12988] = 32'hFFFFFFF1;
    // rom_array[12989] = 32'h0000afe9;
    // rom_array[12990] = 32'h0000aff1;
    // rom_array[12991] = 32'hFFFFFFF1;
    // rom_array[12992] = 32'hFFFFFFF1;
    // rom_array[12993] = 32'h0000aff9;
    // rom_array[12994] = 32'h0000b001;
    // rom_array[12995] = 32'h0000b009;
    // rom_array[12996] = 32'h0000b011;
    // rom_array[12997] = 32'hFFFFFFF0;
    // rom_array[12998] = 32'hFFFFFFF0;
    // rom_array[12999] = 32'hFFFFFFF0;
    // rom_array[13000] = 32'hFFFFFFF0;
    // rom_array[13001] = 32'h0000b019;
    // rom_array[13002] = 32'h0000b021;
    // rom_array[13003] = 32'h0000b029;
    // rom_array[13004] = 32'h0000b031;
    // rom_array[13005] = 32'hFFFFFFF0;
    // rom_array[13006] = 32'hFFFFFFF0;
    // rom_array[13007] = 32'hFFFFFFF0;
    // rom_array[13008] = 32'hFFFFFFF0;
    // rom_array[13009] = 32'h0000b039;
    // rom_array[13010] = 32'h0000b041;
    // rom_array[13011] = 32'h0000b049;
    // rom_array[13012] = 32'h0000b051;
    // rom_array[13013] = 32'hFFFFFFF0;
    // rom_array[13014] = 32'hFFFFFFF0;
    // rom_array[13015] = 32'hFFFFFFF0;
    // rom_array[13016] = 32'hFFFFFFF0;
    // rom_array[13017] = 32'h0000b059;
    // rom_array[13018] = 32'h0000b061;
    // rom_array[13019] = 32'h0000b069;
    // rom_array[13020] = 32'h0000b071;
    // rom_array[13021] = 32'hFFFFFFF0;
    // rom_array[13022] = 32'hFFFFFFF0;
    // rom_array[13023] = 32'hFFFFFFF0;
    // rom_array[13024] = 32'hFFFFFFF0;
    // rom_array[13025] = 32'h0000b079;
    // rom_array[13026] = 32'h0000b081;
    // rom_array[13027] = 32'h0000b089;
    // rom_array[13028] = 32'h0000b091;
    // rom_array[13029] = 32'hFFFFFFF1;
    // rom_array[13030] = 32'hFFFFFFF1;
    // rom_array[13031] = 32'hFFFFFFF1;
    // rom_array[13032] = 32'hFFFFFFF1;
    // rom_array[13033] = 32'h0000b099;
    // rom_array[13034] = 32'h0000b0a1;
    // rom_array[13035] = 32'hFFFFFFF0;
    // rom_array[13036] = 32'hFFFFFFF0;
    // rom_array[13037] = 32'h0000b0a9;
    // rom_array[13038] = 32'h0000b0b1;
    // rom_array[13039] = 32'hFFFFFFF0;
    // rom_array[13040] = 32'hFFFFFFF0;
    // rom_array[13041] = 32'h0000b0b9;
    // rom_array[13042] = 32'h0000b0c1;
    // rom_array[13043] = 32'hFFFFFFF0;
    // rom_array[13044] = 32'hFFFFFFF0;
    // rom_array[13045] = 32'h0000b0c9;
    // rom_array[13046] = 32'h0000b0d1;
    // rom_array[13047] = 32'hFFFFFFF0;
    // rom_array[13048] = 32'hFFFFFFF0;
    // rom_array[13049] = 32'h0000b0d9;
    // rom_array[13050] = 32'h0000b0e1;
    // rom_array[13051] = 32'h0000b0e9;
    // rom_array[13052] = 32'h0000b0f1;
    // rom_array[13053] = 32'hFFFFFFF0;
    // rom_array[13054] = 32'hFFFFFFF0;
    // rom_array[13055] = 32'hFFFFFFF0;
    // rom_array[13056] = 32'hFFFFFFF0;
    // rom_array[13057] = 32'h0000b0f9;
    // rom_array[13058] = 32'h0000b101;
    // rom_array[13059] = 32'hFFFFFFF0;
    // rom_array[13060] = 32'hFFFFFFF0;
    // rom_array[13061] = 32'h0000b109;
    // rom_array[13062] = 32'h0000b111;
    // rom_array[13063] = 32'hFFFFFFF0;
    // rom_array[13064] = 32'hFFFFFFF0;
    // rom_array[13065] = 32'h0000b119;
    // rom_array[13066] = 32'h0000b121;
    // rom_array[13067] = 32'hFFFFFFF0;
    // rom_array[13068] = 32'hFFFFFFF0;
    // rom_array[13069] = 32'h0000b129;
    // rom_array[13070] = 32'h0000b131;
    // rom_array[13071] = 32'hFFFFFFF0;
    // rom_array[13072] = 32'hFFFFFFF0;
    // rom_array[13073] = 32'h0000b139;
    // rom_array[13074] = 32'h0000b141;
    // rom_array[13075] = 32'h0000b149;
    // rom_array[13076] = 32'h0000b151;
    // rom_array[13077] = 32'hFFFFFFF0;
    // rom_array[13078] = 32'hFFFFFFF0;
    // rom_array[13079] = 32'hFFFFFFF0;
    // rom_array[13080] = 32'hFFFFFFF0;
    // rom_array[13081] = 32'h0000b159;
    // rom_array[13082] = 32'h0000b161;
    // rom_array[13083] = 32'h0000b169;
    // rom_array[13084] = 32'h0000b171;
    // rom_array[13085] = 32'hFFFFFFF0;
    // rom_array[13086] = 32'hFFFFFFF0;
    // rom_array[13087] = 32'hFFFFFFF0;
    // rom_array[13088] = 32'hFFFFFFF0;
    // rom_array[13089] = 32'h0000b179;
    // rom_array[13090] = 32'h0000b181;
    // rom_array[13091] = 32'h0000b189;
    // rom_array[13092] = 32'h0000b191;
    // rom_array[13093] = 32'hFFFFFFF0;
    // rom_array[13094] = 32'hFFFFFFF0;
    // rom_array[13095] = 32'hFFFFFFF0;
    // rom_array[13096] = 32'hFFFFFFF0;
    // rom_array[13097] = 32'h0000b199;
    // rom_array[13098] = 32'h0000b1a1;
    // rom_array[13099] = 32'h0000b1a9;
    // rom_array[13100] = 32'h0000b1b1;
    // rom_array[13101] = 32'hFFFFFFF0;
    // rom_array[13102] = 32'hFFFFFFF0;
    // rom_array[13103] = 32'hFFFFFFF0;
    // rom_array[13104] = 32'hFFFFFFF0;
    // rom_array[13105] = 32'h0000b1b9;
    // rom_array[13106] = 32'h0000b1c1;
    // rom_array[13107] = 32'hFFFFFFF0;
    // rom_array[13108] = 32'hFFFFFFF0;
    // rom_array[13109] = 32'h0000b1c9;
    // rom_array[13110] = 32'h0000b1d1;
    // rom_array[13111] = 32'hFFFFFFF0;
    // rom_array[13112] = 32'hFFFFFFF0;
    // rom_array[13113] = 32'h0000b1d9;
    // rom_array[13114] = 32'h0000b1e1;
    // rom_array[13115] = 32'hFFFFFFF0;
    // rom_array[13116] = 32'hFFFFFFF0;
    // rom_array[13117] = 32'h0000b1e9;
    // rom_array[13118] = 32'h0000b1f1;
    // rom_array[13119] = 32'hFFFFFFF0;
    // rom_array[13120] = 32'hFFFFFFF0;
    // rom_array[13121] = 32'h0000b1f9;
    // rom_array[13122] = 32'h0000b201;
    // rom_array[13123] = 32'h0000b209;
    // rom_array[13124] = 32'h0000b211;
    // rom_array[13125] = 32'hFFFFFFF0;
    // rom_array[13126] = 32'hFFFFFFF0;
    // rom_array[13127] = 32'hFFFFFFF0;
    // rom_array[13128] = 32'hFFFFFFF0;
    // rom_array[13129] = 32'h0000b219;
    // rom_array[13130] = 32'h0000b221;
    // rom_array[13131] = 32'hFFFFFFF0;
    // rom_array[13132] = 32'hFFFFFFF0;
    // rom_array[13133] = 32'hFFFFFFF0;
    // rom_array[13134] = 32'hFFFFFFF0;
    // rom_array[13135] = 32'hFFFFFFF0;
    // rom_array[13136] = 32'hFFFFFFF0;
    // rom_array[13137] = 32'h0000b229;
    // rom_array[13138] = 32'h0000b231;
    // rom_array[13139] = 32'h0000b239;
    // rom_array[13140] = 32'h0000b241;
    // rom_array[13141] = 32'hFFFFFFF1;
    // rom_array[13142] = 32'hFFFFFFF1;
    // rom_array[13143] = 32'hFFFFFFF1;
    // rom_array[13144] = 32'hFFFFFFF1;
    // rom_array[13145] = 32'h0000b249;
    // rom_array[13146] = 32'h0000b251;
    // rom_array[13147] = 32'h0000b259;
    // rom_array[13148] = 32'h0000b261;
    // rom_array[13149] = 32'hFFFFFFF1;
    // rom_array[13150] = 32'hFFFFFFF1;
    // rom_array[13151] = 32'hFFFFFFF1;
    // rom_array[13152] = 32'hFFFFFFF1;
    // rom_array[13153] = 32'h0000b269;
    // rom_array[13154] = 32'h0000b271;
    // rom_array[13155] = 32'h0000b279;
    // rom_array[13156] = 32'h0000b281;
    // rom_array[13157] = 32'hFFFFFFF1;
    // rom_array[13158] = 32'hFFFFFFF1;
    // rom_array[13159] = 32'hFFFFFFF1;
    // rom_array[13160] = 32'hFFFFFFF1;
    // rom_array[13161] = 32'h0000b289;
    // rom_array[13162] = 32'h0000b291;
    // rom_array[13163] = 32'h0000b299;
    // rom_array[13164] = 32'h0000b2a1;
    // rom_array[13165] = 32'hFFFFFFF1;
    // rom_array[13166] = 32'hFFFFFFF1;
    // rom_array[13167] = 32'hFFFFFFF1;
    // rom_array[13168] = 32'hFFFFFFF1;
    // rom_array[13169] = 32'h0000b2a9;
    // rom_array[13170] = 32'h0000b2b1;
    // rom_array[13171] = 32'h0000b2b9;
    // rom_array[13172] = 32'h0000b2c1;
    // rom_array[13173] = 32'hFFFFFFF1;
    // rom_array[13174] = 32'hFFFFFFF1;
    // rom_array[13175] = 32'hFFFFFFF1;
    // rom_array[13176] = 32'hFFFFFFF1;
    // rom_array[13177] = 32'h0000b2c9;
    // rom_array[13178] = 32'h0000b2d1;
    // rom_array[13179] = 32'hFFFFFFF0;
    // rom_array[13180] = 32'hFFFFFFF0;
    // rom_array[13181] = 32'h0000b2d9;
    // rom_array[13182] = 32'h0000b2e1;
    // rom_array[13183] = 32'hFFFFFFF0;
    // rom_array[13184] = 32'hFFFFFFF0;
    // rom_array[13185] = 32'h0000b2e9;
    // rom_array[13186] = 32'h0000b2f1;
    // rom_array[13187] = 32'hFFFFFFF0;
    // rom_array[13188] = 32'hFFFFFFF0;
    // rom_array[13189] = 32'h0000b2f9;
    // rom_array[13190] = 32'h0000b301;
    // rom_array[13191] = 32'hFFFFFFF0;
    // rom_array[13192] = 32'hFFFFFFF0;
    // rom_array[13193] = 32'h0000b309;
    // rom_array[13194] = 32'h0000b311;
    // rom_array[13195] = 32'h0000b319;
    // rom_array[13196] = 32'h0000b321;
    // rom_array[13197] = 32'hFFFFFFF0;
    // rom_array[13198] = 32'hFFFFFFF0;
    // rom_array[13199] = 32'hFFFFFFF0;
    // rom_array[13200] = 32'hFFFFFFF0;
    // rom_array[13201] = 32'h0000b329;
    // rom_array[13202] = 32'h0000b331;
    // rom_array[13203] = 32'h0000b339;
    // rom_array[13204] = 32'h0000b341;
    // rom_array[13205] = 32'hFFFFFFF0;
    // rom_array[13206] = 32'hFFFFFFF0;
    // rom_array[13207] = 32'hFFFFFFF0;
    // rom_array[13208] = 32'hFFFFFFF0;
    // rom_array[13209] = 32'h0000b349;
    // rom_array[13210] = 32'h0000b351;
    // rom_array[13211] = 32'h0000b359;
    // rom_array[13212] = 32'h0000b361;
    // rom_array[13213] = 32'hFFFFFFF0;
    // rom_array[13214] = 32'hFFFFFFF0;
    // rom_array[13215] = 32'hFFFFFFF0;
    // rom_array[13216] = 32'hFFFFFFF0;
    // rom_array[13217] = 32'h0000b369;
    // rom_array[13218] = 32'h0000b371;
    // rom_array[13219] = 32'h0000b379;
    // rom_array[13220] = 32'h0000b381;
    // rom_array[13221] = 32'hFFFFFFF0;
    // rom_array[13222] = 32'hFFFFFFF0;
    // rom_array[13223] = 32'hFFFFFFF0;
    // rom_array[13224] = 32'hFFFFFFF0;
    // rom_array[13225] = 32'h0000b389;
    // rom_array[13226] = 32'h0000b391;
    // rom_array[13227] = 32'h0000b399;
    // rom_array[13228] = 32'h0000b3a1;
    // rom_array[13229] = 32'hFFFFFFF0;
    // rom_array[13230] = 32'hFFFFFFF0;
    // rom_array[13231] = 32'hFFFFFFF0;
    // rom_array[13232] = 32'hFFFFFFF0;
    // rom_array[13233] = 32'h0000b3a9;
    // rom_array[13234] = 32'h0000b3b1;
    // rom_array[13235] = 32'hFFFFFFF0;
    // rom_array[13236] = 32'hFFFFFFF0;
    // rom_array[13237] = 32'hFFFFFFF0;
    // rom_array[13238] = 32'hFFFFFFF0;
    // rom_array[13239] = 32'hFFFFFFF0;
    // rom_array[13240] = 32'hFFFFFFF0;
    // rom_array[13241] = 32'hFFFFFFF0;
    // rom_array[13242] = 32'hFFFFFFF0;
    // rom_array[13243] = 32'hFFFFFFF0;
    // rom_array[13244] = 32'hFFFFFFF0;
    // rom_array[13245] = 32'hFFFFFFF0;
    // rom_array[13246] = 32'hFFFFFFF0;
    // rom_array[13247] = 32'hFFFFFFF1;
    // rom_array[13248] = 32'hFFFFFFF1;
    // rom_array[13249] = 32'hFFFFFFF0;
    // rom_array[13250] = 32'hFFFFFFF0;
    // rom_array[13251] = 32'hFFFFFFF0;
    // rom_array[13252] = 32'hFFFFFFF0;
    // rom_array[13253] = 32'hFFFFFFF0;
    // rom_array[13254] = 32'hFFFFFFF0;
    // rom_array[13255] = 32'hFFFFFFF1;
    // rom_array[13256] = 32'hFFFFFFF1;
    // rom_array[13257] = 32'hFFFFFFF0;
    // rom_array[13258] = 32'hFFFFFFF0;
    // rom_array[13259] = 32'hFFFFFFF0;
    // rom_array[13260] = 32'hFFFFFFF0;
    // rom_array[13261] = 32'hFFFFFFF1;
    // rom_array[13262] = 32'hFFFFFFF1;
    // rom_array[13263] = 32'hFFFFFFF1;
    // rom_array[13264] = 32'hFFFFFFF1;
    // rom_array[13265] = 32'hFFFFFFF0;
    // rom_array[13266] = 32'hFFFFFFF0;
    // rom_array[13267] = 32'hFFFFFFF0;
    // rom_array[13268] = 32'hFFFFFFF0;
    // rom_array[13269] = 32'hFFFFFFF1;
    // rom_array[13270] = 32'hFFFFFFF1;
    // rom_array[13271] = 32'hFFFFFFF1;
    // rom_array[13272] = 32'hFFFFFFF1;
    // rom_array[13273] = 32'hFFFFFFF0;
    // rom_array[13274] = 32'hFFFFFFF0;
    // rom_array[13275] = 32'hFFFFFFF0;
    // rom_array[13276] = 32'hFFFFFFF0;
    // rom_array[13277] = 32'hFFFFFFF1;
    // rom_array[13278] = 32'hFFFFFFF1;
    // rom_array[13279] = 32'hFFFFFFF1;
    // rom_array[13280] = 32'hFFFFFFF1;
    // rom_array[13281] = 32'hFFFFFFF0;
    // rom_array[13282] = 32'hFFFFFFF0;
    // rom_array[13283] = 32'hFFFFFFF0;
    // rom_array[13284] = 32'hFFFFFFF0;
    // rom_array[13285] = 32'hFFFFFFF1;
    // rom_array[13286] = 32'hFFFFFFF1;
    // rom_array[13287] = 32'hFFFFFFF1;
    // rom_array[13288] = 32'hFFFFFFF1;
    // rom_array[13289] = 32'hFFFFFFF0;
    // rom_array[13290] = 32'hFFFFFFF0;
    // rom_array[13291] = 32'hFFFFFFF0;
    // rom_array[13292] = 32'hFFFFFFF0;
    // rom_array[13293] = 32'hFFFFFFF1;
    // rom_array[13294] = 32'hFFFFFFF1;
    // rom_array[13295] = 32'hFFFFFFF1;
    // rom_array[13296] = 32'hFFFFFFF1;
    // rom_array[13297] = 32'hFFFFFFF0;
    // rom_array[13298] = 32'hFFFFFFF0;
    // rom_array[13299] = 32'hFFFFFFF0;
    // rom_array[13300] = 32'hFFFFFFF0;
    // rom_array[13301] = 32'hFFFFFFF1;
    // rom_array[13302] = 32'hFFFFFFF1;
    // rom_array[13303] = 32'hFFFFFFF1;
    // rom_array[13304] = 32'hFFFFFFF1;
    // rom_array[13305] = 32'hFFFFFFF0;
    // rom_array[13306] = 32'hFFFFFFF0;
    // rom_array[13307] = 32'hFFFFFFF1;
    // rom_array[13308] = 32'hFFFFFFF1;
    // rom_array[13309] = 32'hFFFFFFF0;
    // rom_array[13310] = 32'hFFFFFFF0;
    // rom_array[13311] = 32'hFFFFFFF1;
    // rom_array[13312] = 32'hFFFFFFF1;
    // rom_array[13313] = 32'hFFFFFFF0;
    // rom_array[13314] = 32'hFFFFFFF0;
    // rom_array[13315] = 32'hFFFFFFF1;
    // rom_array[13316] = 32'hFFFFFFF1;
    // rom_array[13317] = 32'hFFFFFFF0;
    // rom_array[13318] = 32'hFFFFFFF0;
    // rom_array[13319] = 32'hFFFFFFF1;
    // rom_array[13320] = 32'hFFFFFFF1;
    // rom_array[13321] = 32'hFFFFFFF0;
    // rom_array[13322] = 32'hFFFFFFF0;
    // rom_array[13323] = 32'hFFFFFFF1;
    // rom_array[13324] = 32'hFFFFFFF1;
    // rom_array[13325] = 32'hFFFFFFF0;
    // rom_array[13326] = 32'hFFFFFFF0;
    // rom_array[13327] = 32'hFFFFFFF1;
    // rom_array[13328] = 32'hFFFFFFF1;
    // rom_array[13329] = 32'hFFFFFFF0;
    // rom_array[13330] = 32'hFFFFFFF0;
    // rom_array[13331] = 32'hFFFFFFF1;
    // rom_array[13332] = 32'hFFFFFFF1;
    // rom_array[13333] = 32'hFFFFFFF0;
    // rom_array[13334] = 32'hFFFFFFF0;
    // rom_array[13335] = 32'hFFFFFFF1;
    // rom_array[13336] = 32'hFFFFFFF1;
    // rom_array[13337] = 32'hFFFFFFF0;
    // rom_array[13338] = 32'hFFFFFFF0;
    // rom_array[13339] = 32'hFFFFFFF0;
    // rom_array[13340] = 32'hFFFFFFF0;
    // rom_array[13341] = 32'hFFFFFFF1;
    // rom_array[13342] = 32'hFFFFFFF1;
    // rom_array[13343] = 32'hFFFFFFF1;
    // rom_array[13344] = 32'hFFFFFFF1;
    // rom_array[13345] = 32'hFFFFFFF0;
    // rom_array[13346] = 32'hFFFFFFF0;
    // rom_array[13347] = 32'hFFFFFFF0;
    // rom_array[13348] = 32'hFFFFFFF0;
    // rom_array[13349] = 32'hFFFFFFF1;
    // rom_array[13350] = 32'hFFFFFFF1;
    // rom_array[13351] = 32'hFFFFFFF1;
    // rom_array[13352] = 32'hFFFFFFF1;
    // rom_array[13353] = 32'hFFFFFFF1;
    // rom_array[13354] = 32'hFFFFFFF1;
    // rom_array[13355] = 32'hFFFFFFF1;
    // rom_array[13356] = 32'hFFFFFFF1;
    // rom_array[13357] = 32'hFFFFFFF1;
    // rom_array[13358] = 32'hFFFFFFF1;
    // rom_array[13359] = 32'hFFFFFFF1;
    // rom_array[13360] = 32'hFFFFFFF1;
    // rom_array[13361] = 32'hFFFFFFF1;
    // rom_array[13362] = 32'hFFFFFFF1;
    // rom_array[13363] = 32'hFFFFFFF1;
    // rom_array[13364] = 32'hFFFFFFF1;
    // rom_array[13365] = 32'hFFFFFFF1;
    // rom_array[13366] = 32'hFFFFFFF1;
    // rom_array[13367] = 32'hFFFFFFF1;
    // rom_array[13368] = 32'hFFFFFFF1;
    // rom_array[13369] = 32'hFFFFFFF1;
    // rom_array[13370] = 32'hFFFFFFF1;
    // rom_array[13371] = 32'hFFFFFFF1;
    // rom_array[13372] = 32'hFFFFFFF1;
    // rom_array[13373] = 32'hFFFFFFF1;
    // rom_array[13374] = 32'hFFFFFFF1;
    // rom_array[13375] = 32'hFFFFFFF1;
    // rom_array[13376] = 32'hFFFFFFF1;
    // rom_array[13377] = 32'hFFFFFFF1;
    // rom_array[13378] = 32'hFFFFFFF1;
    // rom_array[13379] = 32'hFFFFFFF1;
    // rom_array[13380] = 32'hFFFFFFF1;
    // rom_array[13381] = 32'hFFFFFFF1;
    // rom_array[13382] = 32'hFFFFFFF1;
    // rom_array[13383] = 32'hFFFFFFF1;
    // rom_array[13384] = 32'hFFFFFFF1;
    // rom_array[13385] = 32'hFFFFFFF0;
    // rom_array[13386] = 32'hFFFFFFF0;
    // rom_array[13387] = 32'hFFFFFFF1;
    // rom_array[13388] = 32'hFFFFFFF1;
    // rom_array[13389] = 32'hFFFFFFF0;
    // rom_array[13390] = 32'hFFFFFFF0;
    // rom_array[13391] = 32'hFFFFFFF1;
    // rom_array[13392] = 32'hFFFFFFF1;
    // rom_array[13393] = 32'hFFFFFFF0;
    // rom_array[13394] = 32'hFFFFFFF0;
    // rom_array[13395] = 32'hFFFFFFF1;
    // rom_array[13396] = 32'hFFFFFFF1;
    // rom_array[13397] = 32'hFFFFFFF0;
    // rom_array[13398] = 32'hFFFFFFF0;
    // rom_array[13399] = 32'hFFFFFFF1;
    // rom_array[13400] = 32'hFFFFFFF1;
    // rom_array[13401] = 32'hFFFFFFF0;
    // rom_array[13402] = 32'hFFFFFFF0;
    // rom_array[13403] = 32'hFFFFFFF1;
    // rom_array[13404] = 32'hFFFFFFF1;
    // rom_array[13405] = 32'hFFFFFFF0;
    // rom_array[13406] = 32'hFFFFFFF0;
    // rom_array[13407] = 32'hFFFFFFF1;
    // rom_array[13408] = 32'hFFFFFFF1;
    // rom_array[13409] = 32'hFFFFFFF0;
    // rom_array[13410] = 32'hFFFFFFF0;
    // rom_array[13411] = 32'hFFFFFFF1;
    // rom_array[13412] = 32'hFFFFFFF1;
    // rom_array[13413] = 32'hFFFFFFF0;
    // rom_array[13414] = 32'hFFFFFFF0;
    // rom_array[13415] = 32'hFFFFFFF1;
    // rom_array[13416] = 32'hFFFFFFF1;
    // rom_array[13417] = 32'hFFFFFFF0;
    // rom_array[13418] = 32'hFFFFFFF0;
    // rom_array[13419] = 32'hFFFFFFF1;
    // rom_array[13420] = 32'hFFFFFFF1;
    // rom_array[13421] = 32'hFFFFFFF0;
    // rom_array[13422] = 32'hFFFFFFF0;
    // rom_array[13423] = 32'hFFFFFFF1;
    // rom_array[13424] = 32'hFFFFFFF1;
    // rom_array[13425] = 32'hFFFFFFF0;
    // rom_array[13426] = 32'hFFFFFFF0;
    // rom_array[13427] = 32'hFFFFFFF1;
    // rom_array[13428] = 32'hFFFFFFF1;
    // rom_array[13429] = 32'hFFFFFFF0;
    // rom_array[13430] = 32'hFFFFFFF0;
    // rom_array[13431] = 32'hFFFFFFF1;
    // rom_array[13432] = 32'hFFFFFFF1;
    // rom_array[13433] = 32'hFFFFFFF0;
    // rom_array[13434] = 32'hFFFFFFF0;
    // rom_array[13435] = 32'hFFFFFFF1;
    // rom_array[13436] = 32'hFFFFFFF1;
    // rom_array[13437] = 32'hFFFFFFF0;
    // rom_array[13438] = 32'hFFFFFFF0;
    // rom_array[13439] = 32'hFFFFFFF1;
    // rom_array[13440] = 32'hFFFFFFF1;
    // rom_array[13441] = 32'hFFFFFFF0;
    // rom_array[13442] = 32'hFFFFFFF0;
    // rom_array[13443] = 32'hFFFFFFF1;
    // rom_array[13444] = 32'hFFFFFFF1;
    // rom_array[13445] = 32'hFFFFFFF0;
    // rom_array[13446] = 32'hFFFFFFF0;
    // rom_array[13447] = 32'hFFFFFFF1;
    // rom_array[13448] = 32'hFFFFFFF1;
    // rom_array[13449] = 32'hFFFFFFF0;
    // rom_array[13450] = 32'hFFFFFFF0;
    // rom_array[13451] = 32'hFFFFFFF1;
    // rom_array[13452] = 32'hFFFFFFF1;
    // rom_array[13453] = 32'hFFFFFFF0;
    // rom_array[13454] = 32'hFFFFFFF0;
    // rom_array[13455] = 32'hFFFFFFF1;
    // rom_array[13456] = 32'hFFFFFFF1;
    // rom_array[13457] = 32'hFFFFFFF0;
    // rom_array[13458] = 32'hFFFFFFF0;
    // rom_array[13459] = 32'hFFFFFFF1;
    // rom_array[13460] = 32'hFFFFFFF1;
    // rom_array[13461] = 32'hFFFFFFF0;
    // rom_array[13462] = 32'hFFFFFFF0;
    // rom_array[13463] = 32'hFFFFFFF1;
    // rom_array[13464] = 32'hFFFFFFF1;
    // rom_array[13465] = 32'hFFFFFFF0;
    // rom_array[13466] = 32'hFFFFFFF0;
    // rom_array[13467] = 32'hFFFFFFF1;
    // rom_array[13468] = 32'hFFFFFFF1;
    // rom_array[13469] = 32'hFFFFFFF0;
    // rom_array[13470] = 32'hFFFFFFF0;
    // rom_array[13471] = 32'hFFFFFFF1;
    // rom_array[13472] = 32'hFFFFFFF1;
    // rom_array[13473] = 32'hFFFFFFF0;
    // rom_array[13474] = 32'hFFFFFFF0;
    // rom_array[13475] = 32'hFFFFFFF1;
    // rom_array[13476] = 32'hFFFFFFF1;
    // rom_array[13477] = 32'hFFFFFFF0;
    // rom_array[13478] = 32'hFFFFFFF0;
    // rom_array[13479] = 32'hFFFFFFF1;
    // rom_array[13480] = 32'hFFFFFFF1;
    // rom_array[13481] = 32'hFFFFFFF0;
    // rom_array[13482] = 32'hFFFFFFF0;
    // rom_array[13483] = 32'hFFFFFFF1;
    // rom_array[13484] = 32'hFFFFFFF1;
    // rom_array[13485] = 32'hFFFFFFF0;
    // rom_array[13486] = 32'hFFFFFFF0;
    // rom_array[13487] = 32'hFFFFFFF1;
    // rom_array[13488] = 32'hFFFFFFF1;
    // rom_array[13489] = 32'hFFFFFFF0;
    // rom_array[13490] = 32'hFFFFFFF0;
    // rom_array[13491] = 32'hFFFFFFF1;
    // rom_array[13492] = 32'hFFFFFFF1;
    // rom_array[13493] = 32'hFFFFFFF0;
    // rom_array[13494] = 32'hFFFFFFF0;
    // rom_array[13495] = 32'hFFFFFFF1;
    // rom_array[13496] = 32'hFFFFFFF1;
    // rom_array[13497] = 32'hFFFFFFF0;
    // rom_array[13498] = 32'hFFFFFFF0;
    // rom_array[13499] = 32'hFFFFFFF1;
    // rom_array[13500] = 32'hFFFFFFF1;
    // rom_array[13501] = 32'hFFFFFFF0;
    // rom_array[13502] = 32'hFFFFFFF0;
    // rom_array[13503] = 32'hFFFFFFF1;
    // rom_array[13504] = 32'hFFFFFFF1;
    // rom_array[13505] = 32'hFFFFFFF0;
    // rom_array[13506] = 32'hFFFFFFF0;
    // rom_array[13507] = 32'hFFFFFFF1;
    // rom_array[13508] = 32'hFFFFFFF1;
    // rom_array[13509] = 32'hFFFFFFF0;
    // rom_array[13510] = 32'hFFFFFFF0;
    // rom_array[13511] = 32'hFFFFFFF1;
    // rom_array[13512] = 32'hFFFFFFF1;
    // rom_array[13513] = 32'hFFFFFFF1;
    // rom_array[13514] = 32'hFFFFFFF1;
    // rom_array[13515] = 32'hFFFFFFF1;
    // rom_array[13516] = 32'hFFFFFFF1;
    // rom_array[13517] = 32'hFFFFFFF1;
    // rom_array[13518] = 32'hFFFFFFF1;
    // rom_array[13519] = 32'hFFFFFFF1;
    // rom_array[13520] = 32'hFFFFFFF1;
    // rom_array[13521] = 32'hFFFFFFF1;
    // rom_array[13522] = 32'hFFFFFFF1;
    // rom_array[13523] = 32'hFFFFFFF1;
    // rom_array[13524] = 32'hFFFFFFF1;
    // rom_array[13525] = 32'hFFFFFFF1;
    // rom_array[13526] = 32'hFFFFFFF1;
    // rom_array[13527] = 32'hFFFFFFF1;
    // rom_array[13528] = 32'hFFFFFFF1;
    // rom_array[13529] = 32'hFFFFFFF1;
    // rom_array[13530] = 32'hFFFFFFF1;
    // rom_array[13531] = 32'hFFFFFFF1;
    // rom_array[13532] = 32'hFFFFFFF1;
    // rom_array[13533] = 32'hFFFFFFF1;
    // rom_array[13534] = 32'hFFFFFFF1;
    // rom_array[13535] = 32'hFFFFFFF1;
    // rom_array[13536] = 32'hFFFFFFF1;
    // rom_array[13537] = 32'hFFFFFFF1;
    // rom_array[13538] = 32'hFFFFFFF1;
    // rom_array[13539] = 32'hFFFFFFF1;
    // rom_array[13540] = 32'hFFFFFFF1;
    // rom_array[13541] = 32'hFFFFFFF1;
    // rom_array[13542] = 32'hFFFFFFF1;
    // rom_array[13543] = 32'hFFFFFFF1;
    // rom_array[13544] = 32'hFFFFFFF1;
    // rom_array[13545] = 32'hFFFFFFF1;
    // rom_array[13546] = 32'hFFFFFFF1;
    // rom_array[13547] = 32'hFFFFFFF1;
    // rom_array[13548] = 32'hFFFFFFF1;
    // rom_array[13549] = 32'hFFFFFFF1;
    // rom_array[13550] = 32'hFFFFFFF1;
    // rom_array[13551] = 32'hFFFFFFF1;
    // rom_array[13552] = 32'hFFFFFFF1;
    // rom_array[13553] = 32'hFFFFFFF1;
    // rom_array[13554] = 32'hFFFFFFF1;
    // rom_array[13555] = 32'hFFFFFFF1;
    // rom_array[13556] = 32'hFFFFFFF1;
    // rom_array[13557] = 32'hFFFFFFF1;
    // rom_array[13558] = 32'hFFFFFFF1;
    // rom_array[13559] = 32'hFFFFFFF1;
    // rom_array[13560] = 32'hFFFFFFF1;
    // rom_array[13561] = 32'hFFFFFFF0;
    // rom_array[13562] = 32'hFFFFFFF0;
    // rom_array[13563] = 32'hFFFFFFF0;
    // rom_array[13564] = 32'hFFFFFFF0;
    // rom_array[13565] = 32'hFFFFFFF1;
    // rom_array[13566] = 32'hFFFFFFF1;
    // rom_array[13567] = 32'hFFFFFFF1;
    // rom_array[13568] = 32'hFFFFFFF1;
    // rom_array[13569] = 32'hFFFFFFF0;
    // rom_array[13570] = 32'hFFFFFFF0;
    // rom_array[13571] = 32'hFFFFFFF0;
    // rom_array[13572] = 32'hFFFFFFF0;
    // rom_array[13573] = 32'hFFFFFFF1;
    // rom_array[13574] = 32'hFFFFFFF1;
    // rom_array[13575] = 32'hFFFFFFF1;
    // rom_array[13576] = 32'hFFFFFFF1;
    // rom_array[13577] = 32'hFFFFFFF1;
    // rom_array[13578] = 32'hFFFFFFF1;
    // rom_array[13579] = 32'hFFFFFFF1;
    // rom_array[13580] = 32'hFFFFFFF1;
    // rom_array[13581] = 32'hFFFFFFF1;
    // rom_array[13582] = 32'hFFFFFFF1;
    // rom_array[13583] = 32'hFFFFFFF1;
    // rom_array[13584] = 32'hFFFFFFF1;
    // rom_array[13585] = 32'hFFFFFFF1;
    // rom_array[13586] = 32'hFFFFFFF1;
    // rom_array[13587] = 32'hFFFFFFF1;
    // rom_array[13588] = 32'hFFFFFFF1;
    // rom_array[13589] = 32'hFFFFFFF1;
    // rom_array[13590] = 32'hFFFFFFF1;
    // rom_array[13591] = 32'hFFFFFFF1;
    // rom_array[13592] = 32'hFFFFFFF1;
    // rom_array[13593] = 32'hFFFFFFF0;
    // rom_array[13594] = 32'hFFFFFFF0;
    // rom_array[13595] = 32'hFFFFFFF0;
    // rom_array[13596] = 32'hFFFFFFF0;
    // rom_array[13597] = 32'hFFFFFFF1;
    // rom_array[13598] = 32'hFFFFFFF1;
    // rom_array[13599] = 32'hFFFFFFF1;
    // rom_array[13600] = 32'hFFFFFFF1;
    // rom_array[13601] = 32'hFFFFFFF0;
    // rom_array[13602] = 32'hFFFFFFF0;
    // rom_array[13603] = 32'hFFFFFFF0;
    // rom_array[13604] = 32'hFFFFFFF0;
    // rom_array[13605] = 32'hFFFFFFF1;
    // rom_array[13606] = 32'hFFFFFFF1;
    // rom_array[13607] = 32'hFFFFFFF1;
    // rom_array[13608] = 32'hFFFFFFF1;
    // rom_array[13609] = 32'hFFFFFFF0;
    // rom_array[13610] = 32'hFFFFFFF0;
    // rom_array[13611] = 32'hFFFFFFF0;
    // rom_array[13612] = 32'hFFFFFFF0;
    // rom_array[13613] = 32'hFFFFFFF1;
    // rom_array[13614] = 32'hFFFFFFF1;
    // rom_array[13615] = 32'hFFFFFFF1;
    // rom_array[13616] = 32'hFFFFFFF1;
    // rom_array[13617] = 32'hFFFFFFF0;
    // rom_array[13618] = 32'hFFFFFFF0;
    // rom_array[13619] = 32'hFFFFFFF0;
    // rom_array[13620] = 32'hFFFFFFF0;
    // rom_array[13621] = 32'hFFFFFFF1;
    // rom_array[13622] = 32'hFFFFFFF1;
    // rom_array[13623] = 32'hFFFFFFF1;
    // rom_array[13624] = 32'hFFFFFFF1;
    // rom_array[13625] = 32'hFFFFFFF0;
    // rom_array[13626] = 32'hFFFFFFF0;
    // rom_array[13627] = 32'hFFFFFFF0;
    // rom_array[13628] = 32'hFFFFFFF0;
    // rom_array[13629] = 32'hFFFFFFF1;
    // rom_array[13630] = 32'hFFFFFFF1;
    // rom_array[13631] = 32'hFFFFFFF1;
    // rom_array[13632] = 32'hFFFFFFF1;
    // rom_array[13633] = 32'hFFFFFFF0;
    // rom_array[13634] = 32'hFFFFFFF0;
    // rom_array[13635] = 32'hFFFFFFF0;
    // rom_array[13636] = 32'hFFFFFFF0;
    // rom_array[13637] = 32'hFFFFFFF1;
    // rom_array[13638] = 32'hFFFFFFF1;
    // rom_array[13639] = 32'hFFFFFFF1;
    // rom_array[13640] = 32'hFFFFFFF1;
    // rom_array[13641] = 32'hFFFFFFF0;
    // rom_array[13642] = 32'hFFFFFFF0;
    // rom_array[13643] = 32'hFFFFFFF0;
    // rom_array[13644] = 32'hFFFFFFF0;
    // rom_array[13645] = 32'hFFFFFFF1;
    // rom_array[13646] = 32'hFFFFFFF1;
    // rom_array[13647] = 32'hFFFFFFF1;
    // rom_array[13648] = 32'hFFFFFFF1;
    // rom_array[13649] = 32'hFFFFFFF0;
    // rom_array[13650] = 32'hFFFFFFF0;
    // rom_array[13651] = 32'hFFFFFFF0;
    // rom_array[13652] = 32'hFFFFFFF0;
    // rom_array[13653] = 32'hFFFFFFF1;
    // rom_array[13654] = 32'hFFFFFFF1;
    // rom_array[13655] = 32'hFFFFFFF1;
    // rom_array[13656] = 32'hFFFFFFF1;
    // rom_array[13657] = 32'hFFFFFFF0;
    // rom_array[13658] = 32'hFFFFFFF0;
    // rom_array[13659] = 32'hFFFFFFF0;
    // rom_array[13660] = 32'hFFFFFFF0;
    // rom_array[13661] = 32'hFFFFFFF1;
    // rom_array[13662] = 32'hFFFFFFF1;
    // rom_array[13663] = 32'hFFFFFFF1;
    // rom_array[13664] = 32'hFFFFFFF1;
    // rom_array[13665] = 32'hFFFFFFF0;
    // rom_array[13666] = 32'hFFFFFFF0;
    // rom_array[13667] = 32'hFFFFFFF0;
    // rom_array[13668] = 32'hFFFFFFF0;
    // rom_array[13669] = 32'hFFFFFFF1;
    // rom_array[13670] = 32'hFFFFFFF1;
    // rom_array[13671] = 32'hFFFFFFF1;
    // rom_array[13672] = 32'hFFFFFFF1;
    // rom_array[13673] = 32'hFFFFFFF0;
    // rom_array[13674] = 32'hFFFFFFF0;
    // rom_array[13675] = 32'hFFFFFFF0;
    // rom_array[13676] = 32'hFFFFFFF0;
    // rom_array[13677] = 32'hFFFFFFF1;
    // rom_array[13678] = 32'hFFFFFFF1;
    // rom_array[13679] = 32'hFFFFFFF1;
    // rom_array[13680] = 32'hFFFFFFF1;
    // rom_array[13681] = 32'hFFFFFFF0;
    // rom_array[13682] = 32'hFFFFFFF0;
    // rom_array[13683] = 32'hFFFFFFF0;
    // rom_array[13684] = 32'hFFFFFFF0;
    // rom_array[13685] = 32'hFFFFFFF1;
    // rom_array[13686] = 32'hFFFFFFF1;
    // rom_array[13687] = 32'hFFFFFFF1;
    // rom_array[13688] = 32'hFFFFFFF1;
    // rom_array[13689] = 32'hFFFFFFF1;
    // rom_array[13690] = 32'hFFFFFFF1;
    // rom_array[13691] = 32'hFFFFFFF1;
    // rom_array[13692] = 32'hFFFFFFF1;
    // rom_array[13693] = 32'hFFFFFFF1;
    // rom_array[13694] = 32'hFFFFFFF1;
    // rom_array[13695] = 32'hFFFFFFF1;
    // rom_array[13696] = 32'hFFFFFFF1;
    // rom_array[13697] = 32'hFFFFFFF1;
    // rom_array[13698] = 32'hFFFFFFF1;
    // rom_array[13699] = 32'hFFFFFFF1;
    // rom_array[13700] = 32'hFFFFFFF1;
    // rom_array[13701] = 32'hFFFFFFF1;
    // rom_array[13702] = 32'hFFFFFFF1;
    // rom_array[13703] = 32'hFFFFFFF1;
    // rom_array[13704] = 32'hFFFFFFF1;
    // rom_array[13705] = 32'hFFFFFFF1;
    // rom_array[13706] = 32'hFFFFFFF1;
    // rom_array[13707] = 32'hFFFFFFF1;
    // rom_array[13708] = 32'hFFFFFFF1;
    // rom_array[13709] = 32'hFFFFFFF1;
    // rom_array[13710] = 32'hFFFFFFF1;
    // rom_array[13711] = 32'hFFFFFFF1;
    // rom_array[13712] = 32'hFFFFFFF1;
    // rom_array[13713] = 32'hFFFFFFF1;
    // rom_array[13714] = 32'hFFFFFFF1;
    // rom_array[13715] = 32'hFFFFFFF1;
    // rom_array[13716] = 32'hFFFFFFF1;
    // rom_array[13717] = 32'hFFFFFFF1;
    // rom_array[13718] = 32'hFFFFFFF1;
    // rom_array[13719] = 32'hFFFFFFF1;
    // rom_array[13720] = 32'hFFFFFFF1;
    // rom_array[13721] = 32'hFFFFFFF1;
    // rom_array[13722] = 32'hFFFFFFF1;
    // rom_array[13723] = 32'hFFFFFFF1;
    // rom_array[13724] = 32'hFFFFFFF1;
    // rom_array[13725] = 32'hFFFFFFF1;
    // rom_array[13726] = 32'hFFFFFFF1;
    // rom_array[13727] = 32'hFFFFFFF1;
    // rom_array[13728] = 32'hFFFFFFF1;
    // rom_array[13729] = 32'hFFFFFFF1;
    // rom_array[13730] = 32'hFFFFFFF1;
    // rom_array[13731] = 32'hFFFFFFF1;
    // rom_array[13732] = 32'hFFFFFFF1;
    // rom_array[13733] = 32'hFFFFFFF1;
    // rom_array[13734] = 32'hFFFFFFF1;
    // rom_array[13735] = 32'hFFFFFFF1;
    // rom_array[13736] = 32'hFFFFFFF1;
    // rom_array[13737] = 32'hFFFFFFF1;
    // rom_array[13738] = 32'hFFFFFFF1;
    // rom_array[13739] = 32'hFFFFFFF1;
    // rom_array[13740] = 32'hFFFFFFF1;
    // rom_array[13741] = 32'hFFFFFFF0;
    // rom_array[13742] = 32'hFFFFFFF0;
    // rom_array[13743] = 32'hFFFFFFF0;
    // rom_array[13744] = 32'hFFFFFFF0;
    // rom_array[13745] = 32'hFFFFFFF1;
    // rom_array[13746] = 32'hFFFFFFF1;
    // rom_array[13747] = 32'hFFFFFFF1;
    // rom_array[13748] = 32'hFFFFFFF1;
    // rom_array[13749] = 32'hFFFFFFF0;
    // rom_array[13750] = 32'hFFFFFFF0;
    // rom_array[13751] = 32'hFFFFFFF0;
    // rom_array[13752] = 32'hFFFFFFF0;
    // rom_array[13753] = 32'hFFFFFFF1;
    // rom_array[13754] = 32'hFFFFFFF1;
    // rom_array[13755] = 32'hFFFFFFF1;
    // rom_array[13756] = 32'hFFFFFFF1;
    // rom_array[13757] = 32'hFFFFFFF1;
    // rom_array[13758] = 32'hFFFFFFF1;
    // rom_array[13759] = 32'hFFFFFFF1;
    // rom_array[13760] = 32'hFFFFFFF1;
    // rom_array[13761] = 32'hFFFFFFF1;
    // rom_array[13762] = 32'hFFFFFFF1;
    // rom_array[13763] = 32'hFFFFFFF1;
    // rom_array[13764] = 32'hFFFFFFF1;
    // rom_array[13765] = 32'hFFFFFFF1;
    // rom_array[13766] = 32'hFFFFFFF1;
    // rom_array[13767] = 32'hFFFFFFF1;
    // rom_array[13768] = 32'hFFFFFFF1;
    // rom_array[13769] = 32'hFFFFFFF1;
    // rom_array[13770] = 32'hFFFFFFF1;
    // rom_array[13771] = 32'hFFFFFFF1;
    // rom_array[13772] = 32'hFFFFFFF1;
    // rom_array[13773] = 32'hFFFFFFF0;
    // rom_array[13774] = 32'hFFFFFFF0;
    // rom_array[13775] = 32'hFFFFFFF0;
    // rom_array[13776] = 32'hFFFFFFF0;
    // rom_array[13777] = 32'hFFFFFFF1;
    // rom_array[13778] = 32'hFFFFFFF1;
    // rom_array[13779] = 32'hFFFFFFF1;
    // rom_array[13780] = 32'hFFFFFFF1;
    // rom_array[13781] = 32'hFFFFFFF0;
    // rom_array[13782] = 32'hFFFFFFF0;
    // rom_array[13783] = 32'hFFFFFFF0;
    // rom_array[13784] = 32'hFFFFFFF0;
    // rom_array[13785] = 32'hFFFFFFF1;
    // rom_array[13786] = 32'hFFFFFFF1;
    // rom_array[13787] = 32'hFFFFFFF1;
    // rom_array[13788] = 32'hFFFFFFF1;
    // rom_array[13789] = 32'hFFFFFFF0;
    // rom_array[13790] = 32'hFFFFFFF0;
    // rom_array[13791] = 32'hFFFFFFF0;
    // rom_array[13792] = 32'hFFFFFFF0;
    // rom_array[13793] = 32'hFFFFFFF1;
    // rom_array[13794] = 32'hFFFFFFF1;
    // rom_array[13795] = 32'hFFFFFFF1;
    // rom_array[13796] = 32'hFFFFFFF1;
    // rom_array[13797] = 32'hFFFFFFF0;
    // rom_array[13798] = 32'hFFFFFFF0;
    // rom_array[13799] = 32'hFFFFFFF0;
    // rom_array[13800] = 32'hFFFFFFF0;
    // rom_array[13801] = 32'hFFFFFFF1;
    // rom_array[13802] = 32'hFFFFFFF1;
    // rom_array[13803] = 32'hFFFFFFF1;
    // rom_array[13804] = 32'hFFFFFFF1;
    // rom_array[13805] = 32'hFFFFFFF0;
    // rom_array[13806] = 32'hFFFFFFF0;
    // rom_array[13807] = 32'hFFFFFFF0;
    // rom_array[13808] = 32'hFFFFFFF0;
    // rom_array[13809] = 32'hFFFFFFF1;
    // rom_array[13810] = 32'hFFFFFFF1;
    // rom_array[13811] = 32'hFFFFFFF1;
    // rom_array[13812] = 32'hFFFFFFF1;
    // rom_array[13813] = 32'hFFFFFFF0;
    // rom_array[13814] = 32'hFFFFFFF0;
    // rom_array[13815] = 32'hFFFFFFF0;
    // rom_array[13816] = 32'hFFFFFFF0;
    // rom_array[13817] = 32'hFFFFFFF1;
    // rom_array[13818] = 32'hFFFFFFF1;
    // rom_array[13819] = 32'hFFFFFFF1;
    // rom_array[13820] = 32'hFFFFFFF1;
    // rom_array[13821] = 32'hFFFFFFF0;
    // rom_array[13822] = 32'hFFFFFFF0;
    // rom_array[13823] = 32'hFFFFFFF0;
    // rom_array[13824] = 32'hFFFFFFF0;
    // rom_array[13825] = 32'hFFFFFFF1;
    // rom_array[13826] = 32'hFFFFFFF1;
    // rom_array[13827] = 32'hFFFFFFF1;
    // rom_array[13828] = 32'hFFFFFFF1;
    // rom_array[13829] = 32'hFFFFFFF0;
    // rom_array[13830] = 32'hFFFFFFF0;
    // rom_array[13831] = 32'hFFFFFFF0;
    // rom_array[13832] = 32'hFFFFFFF0;
    // rom_array[13833] = 32'hFFFFFFF1;
    // rom_array[13834] = 32'hFFFFFFF1;
    // rom_array[13835] = 32'hFFFFFFF1;
    // rom_array[13836] = 32'hFFFFFFF1;
    // rom_array[13837] = 32'hFFFFFFF0;
    // rom_array[13838] = 32'hFFFFFFF0;
    // rom_array[13839] = 32'hFFFFFFF0;
    // rom_array[13840] = 32'hFFFFFFF0;
    // rom_array[13841] = 32'hFFFFFFF1;
    // rom_array[13842] = 32'hFFFFFFF1;
    // rom_array[13843] = 32'hFFFFFFF1;
    // rom_array[13844] = 32'hFFFFFFF1;
    // rom_array[13845] = 32'hFFFFFFF0;
    // rom_array[13846] = 32'hFFFFFFF0;
    // rom_array[13847] = 32'hFFFFFFF0;
    // rom_array[13848] = 32'hFFFFFFF0;
    // rom_array[13849] = 32'hFFFFFFF1;
    // rom_array[13850] = 32'hFFFFFFF1;
    // rom_array[13851] = 32'hFFFFFFF1;
    // rom_array[13852] = 32'hFFFFFFF1;
    // rom_array[13853] = 32'hFFFFFFF0;
    // rom_array[13854] = 32'hFFFFFFF0;
    // rom_array[13855] = 32'hFFFFFFF0;
    // rom_array[13856] = 32'hFFFFFFF0;
    // rom_array[13857] = 32'hFFFFFFF1;
    // rom_array[13858] = 32'hFFFFFFF1;
    // rom_array[13859] = 32'hFFFFFFF1;
    // rom_array[13860] = 32'hFFFFFFF1;
    // rom_array[13861] = 32'hFFFFFFF0;
    // rom_array[13862] = 32'hFFFFFFF0;
    // rom_array[13863] = 32'hFFFFFFF0;
    // rom_array[13864] = 32'hFFFFFFF0;
    // rom_array[13865] = 32'hFFFFFFF0;
    // rom_array[13866] = 32'hFFFFFFF0;
    // rom_array[13867] = 32'hFFFFFFF1;
    // rom_array[13868] = 32'hFFFFFFF1;
    // rom_array[13869] = 32'hFFFFFFF0;
    // rom_array[13870] = 32'hFFFFFFF0;
    // rom_array[13871] = 32'hFFFFFFF1;
    // rom_array[13872] = 32'hFFFFFFF1;
    // rom_array[13873] = 32'hFFFFFFF0;
    // rom_array[13874] = 32'hFFFFFFF0;
    // rom_array[13875] = 32'hFFFFFFF1;
    // rom_array[13876] = 32'hFFFFFFF1;
    // rom_array[13877] = 32'hFFFFFFF0;
    // rom_array[13878] = 32'hFFFFFFF0;
    // rom_array[13879] = 32'hFFFFFFF1;
    // rom_array[13880] = 32'hFFFFFFF1;
    // rom_array[13881] = 32'hFFFFFFF0;
    // rom_array[13882] = 32'hFFFFFFF0;
    // rom_array[13883] = 32'hFFFFFFF1;
    // rom_array[13884] = 32'hFFFFFFF1;
    // rom_array[13885] = 32'hFFFFFFF0;
    // rom_array[13886] = 32'hFFFFFFF0;
    // rom_array[13887] = 32'hFFFFFFF1;
    // rom_array[13888] = 32'hFFFFFFF1;
    // rom_array[13889] = 32'hFFFFFFF0;
    // rom_array[13890] = 32'hFFFFFFF0;
    // rom_array[13891] = 32'hFFFFFFF1;
    // rom_array[13892] = 32'hFFFFFFF1;
    // rom_array[13893] = 32'hFFFFFFF0;
    // rom_array[13894] = 32'hFFFFFFF0;
    // rom_array[13895] = 32'hFFFFFFF1;
    // rom_array[13896] = 32'hFFFFFFF1;
    // rom_array[13897] = 32'hFFFFFFF0;
    // rom_array[13898] = 32'hFFFFFFF0;
    // rom_array[13899] = 32'hFFFFFFF1;
    // rom_array[13900] = 32'hFFFFFFF1;
    // rom_array[13901] = 32'hFFFFFFF0;
    // rom_array[13902] = 32'hFFFFFFF0;
    // rom_array[13903] = 32'hFFFFFFF1;
    // rom_array[13904] = 32'hFFFFFFF1;
    // rom_array[13905] = 32'hFFFFFFF0;
    // rom_array[13906] = 32'hFFFFFFF0;
    // rom_array[13907] = 32'hFFFFFFF1;
    // rom_array[13908] = 32'hFFFFFFF1;
    // rom_array[13909] = 32'hFFFFFFF0;
    // rom_array[13910] = 32'hFFFFFFF0;
    // rom_array[13911] = 32'hFFFFFFF1;
    // rom_array[13912] = 32'hFFFFFFF1;
    // rom_array[13913] = 32'hFFFFFFF0;
    // rom_array[13914] = 32'hFFFFFFF0;
    // rom_array[13915] = 32'hFFFFFFF1;
    // rom_array[13916] = 32'hFFFFFFF1;
    // rom_array[13917] = 32'hFFFFFFF0;
    // rom_array[13918] = 32'hFFFFFFF0;
    // rom_array[13919] = 32'hFFFFFFF0;
    // rom_array[13920] = 32'hFFFFFFF0;
    // rom_array[13921] = 32'hFFFFFFF0;
    // rom_array[13922] = 32'hFFFFFFF0;
    // rom_array[13923] = 32'hFFFFFFF1;
    // rom_array[13924] = 32'hFFFFFFF1;
    // rom_array[13925] = 32'hFFFFFFF0;
    // rom_array[13926] = 32'hFFFFFFF0;
    // rom_array[13927] = 32'hFFFFFFF0;
    // rom_array[13928] = 32'hFFFFFFF0;
    // rom_array[13929] = 32'hFFFFFFF1;
    // rom_array[13930] = 32'hFFFFFFF1;
    // rom_array[13931] = 32'hFFFFFFF1;
    // rom_array[13932] = 32'hFFFFFFF1;
    // rom_array[13933] = 32'hFFFFFFF0;
    // rom_array[13934] = 32'hFFFFFFF0;
    // rom_array[13935] = 32'hFFFFFFF0;
    // rom_array[13936] = 32'hFFFFFFF0;
    // rom_array[13937] = 32'hFFFFFFF1;
    // rom_array[13938] = 32'hFFFFFFF1;
    // rom_array[13939] = 32'hFFFFFFF1;
    // rom_array[13940] = 32'hFFFFFFF1;
    // rom_array[13941] = 32'hFFFFFFF0;
    // rom_array[13942] = 32'hFFFFFFF0;
    // rom_array[13943] = 32'hFFFFFFF0;
    // rom_array[13944] = 32'hFFFFFFF0;
    // rom_array[13945] = 32'hFFFFFFF1;
    // rom_array[13946] = 32'hFFFFFFF1;
    // rom_array[13947] = 32'hFFFFFFF1;
    // rom_array[13948] = 32'hFFFFFFF1;
    // rom_array[13949] = 32'hFFFFFFF0;
    // rom_array[13950] = 32'hFFFFFFF0;
    // rom_array[13951] = 32'hFFFFFFF0;
    // rom_array[13952] = 32'hFFFFFFF0;
    // rom_array[13953] = 32'hFFFFFFF1;
    // rom_array[13954] = 32'hFFFFFFF1;
    // rom_array[13955] = 32'hFFFFFFF1;
    // rom_array[13956] = 32'hFFFFFFF1;
    // rom_array[13957] = 32'hFFFFFFF0;
    // rom_array[13958] = 32'hFFFFFFF0;
    // rom_array[13959] = 32'hFFFFFFF0;
    // rom_array[13960] = 32'hFFFFFFF0;
    // rom_array[13961] = 32'hFFFFFFF1;
    // rom_array[13962] = 32'hFFFFFFF1;
    // rom_array[13963] = 32'hFFFFFFF1;
    // rom_array[13964] = 32'hFFFFFFF1;
    // rom_array[13965] = 32'hFFFFFFF0;
    // rom_array[13966] = 32'hFFFFFFF0;
    // rom_array[13967] = 32'hFFFFFFF0;
    // rom_array[13968] = 32'hFFFFFFF0;
    // rom_array[13969] = 32'hFFFFFFF1;
    // rom_array[13970] = 32'hFFFFFFF1;
    // rom_array[13971] = 32'hFFFFFFF1;
    // rom_array[13972] = 32'hFFFFFFF1;
    // rom_array[13973] = 32'hFFFFFFF0;
    // rom_array[13974] = 32'hFFFFFFF0;
    // rom_array[13975] = 32'hFFFFFFF0;
    // rom_array[13976] = 32'hFFFFFFF0;
    // rom_array[13977] = 32'hFFFFFFF1;
    // rom_array[13978] = 32'hFFFFFFF1;
    // rom_array[13979] = 32'hFFFFFFF1;
    // rom_array[13980] = 32'hFFFFFFF1;
    // rom_array[13981] = 32'hFFFFFFF1;
    // rom_array[13982] = 32'hFFFFFFF1;
    // rom_array[13983] = 32'hFFFFFFF1;
    // rom_array[13984] = 32'hFFFFFFF1;
    // rom_array[13985] = 32'hFFFFFFF1;
    // rom_array[13986] = 32'hFFFFFFF1;
    // rom_array[13987] = 32'hFFFFFFF1;
    // rom_array[13988] = 32'hFFFFFFF1;
    // rom_array[13989] = 32'hFFFFFFF1;
    // rom_array[13990] = 32'hFFFFFFF1;
    // rom_array[13991] = 32'hFFFFFFF1;
    // rom_array[13992] = 32'hFFFFFFF1;
    // rom_array[13993] = 32'hFFFFFFF1;
    // rom_array[13994] = 32'hFFFFFFF1;
    // rom_array[13995] = 32'hFFFFFFF1;
    // rom_array[13996] = 32'hFFFFFFF1;
    // rom_array[13997] = 32'hFFFFFFF1;
    // rom_array[13998] = 32'hFFFFFFF1;
    // rom_array[13999] = 32'hFFFFFFF1;
    // rom_array[14000] = 32'hFFFFFFF1;
    // rom_array[14001] = 32'hFFFFFFF1;
    // rom_array[14002] = 32'hFFFFFFF1;
    // rom_array[14003] = 32'hFFFFFFF1;
    // rom_array[14004] = 32'hFFFFFFF1;
    // rom_array[14005] = 32'hFFFFFFF1;
    // rom_array[14006] = 32'hFFFFFFF1;
    // rom_array[14007] = 32'hFFFFFFF1;
    // rom_array[14008] = 32'hFFFFFFF1;
    // rom_array[14009] = 32'hFFFFFFF1;
    // rom_array[14010] = 32'hFFFFFFF1;
    // rom_array[14011] = 32'hFFFFFFF1;
    // rom_array[14012] = 32'hFFFFFFF1;
    // rom_array[14013] = 32'hFFFFFFF1;
    // rom_array[14014] = 32'hFFFFFFF1;
    // rom_array[14015] = 32'hFFFFFFF1;
    // rom_array[14016] = 32'hFFFFFFF1;
    // rom_array[14017] = 32'hFFFFFFF1;
    // rom_array[14018] = 32'hFFFFFFF1;
    // rom_array[14019] = 32'hFFFFFFF1;
    // rom_array[14020] = 32'hFFFFFFF1;
    // rom_array[14021] = 32'hFFFFFFF1;
    // rom_array[14022] = 32'hFFFFFFF1;
    // rom_array[14023] = 32'hFFFFFFF1;
    // rom_array[14024] = 32'hFFFFFFF1;
    // rom_array[14025] = 32'hFFFFFFF1;
    // rom_array[14026] = 32'hFFFFFFF1;
    // rom_array[14027] = 32'hFFFFFFF1;
    // rom_array[14028] = 32'hFFFFFFF1;
    // rom_array[14029] = 32'hFFFFFFF0;
    // rom_array[14030] = 32'hFFFFFFF0;
    // rom_array[14031] = 32'hFFFFFFF0;
    // rom_array[14032] = 32'hFFFFFFF0;
    // rom_array[14033] = 32'hFFFFFFF1;
    // rom_array[14034] = 32'hFFFFFFF1;
    // rom_array[14035] = 32'hFFFFFFF1;
    // rom_array[14036] = 32'hFFFFFFF1;
    // rom_array[14037] = 32'hFFFFFFF0;
    // rom_array[14038] = 32'hFFFFFFF0;
    // rom_array[14039] = 32'hFFFFFFF0;
    // rom_array[14040] = 32'hFFFFFFF0;
    // rom_array[14041] = 32'hFFFFFFF0;
    // rom_array[14042] = 32'hFFFFFFF0;
    // rom_array[14043] = 32'hFFFFFFF0;
    // rom_array[14044] = 32'hFFFFFFF0;
    // rom_array[14045] = 32'hFFFFFFF0;
    // rom_array[14046] = 32'hFFFFFFF0;
    // rom_array[14047] = 32'hFFFFFFF1;
    // rom_array[14048] = 32'hFFFFFFF1;
    // rom_array[14049] = 32'hFFFFFFF0;
    // rom_array[14050] = 32'hFFFFFFF0;
    // rom_array[14051] = 32'hFFFFFFF0;
    // rom_array[14052] = 32'hFFFFFFF0;
    // rom_array[14053] = 32'hFFFFFFF0;
    // rom_array[14054] = 32'hFFFFFFF0;
    // rom_array[14055] = 32'hFFFFFFF1;
    // rom_array[14056] = 32'hFFFFFFF1;
    // rom_array[14057] = 32'hFFFFFFF0;
    // rom_array[14058] = 32'hFFFFFFF0;
    // rom_array[14059] = 32'hFFFFFFF0;
    // rom_array[14060] = 32'hFFFFFFF0;
    // rom_array[14061] = 32'hFFFFFFF1;
    // rom_array[14062] = 32'hFFFFFFF1;
    // rom_array[14063] = 32'hFFFFFFF1;
    // rom_array[14064] = 32'hFFFFFFF1;
    // rom_array[14065] = 32'hFFFFFFF0;
    // rom_array[14066] = 32'hFFFFFFF0;
    // rom_array[14067] = 32'hFFFFFFF0;
    // rom_array[14068] = 32'hFFFFFFF0;
    // rom_array[14069] = 32'hFFFFFFF1;
    // rom_array[14070] = 32'hFFFFFFF1;
    // rom_array[14071] = 32'hFFFFFFF1;
    // rom_array[14072] = 32'hFFFFFFF1;
    // rom_array[14073] = 32'hFFFFFFF0;
    // rom_array[14074] = 32'hFFFFFFF0;
    // rom_array[14075] = 32'hFFFFFFF1;
    // rom_array[14076] = 32'hFFFFFFF1;
    // rom_array[14077] = 32'hFFFFFFF0;
    // rom_array[14078] = 32'hFFFFFFF0;
    // rom_array[14079] = 32'hFFFFFFF1;
    // rom_array[14080] = 32'hFFFFFFF1;
    // rom_array[14081] = 32'hFFFFFFF0;
    // rom_array[14082] = 32'hFFFFFFF0;
    // rom_array[14083] = 32'hFFFFFFF1;
    // rom_array[14084] = 32'hFFFFFFF1;
    // rom_array[14085] = 32'hFFFFFFF0;
    // rom_array[14086] = 32'hFFFFFFF0;
    // rom_array[14087] = 32'hFFFFFFF1;
    // rom_array[14088] = 32'hFFFFFFF1;
    // rom_array[14089] = 32'hFFFFFFF0;
    // rom_array[14090] = 32'hFFFFFFF0;
    // rom_array[14091] = 32'hFFFFFFF0;
    // rom_array[14092] = 32'hFFFFFFF0;
    // rom_array[14093] = 32'hFFFFFFF1;
    // rom_array[14094] = 32'hFFFFFFF1;
    // rom_array[14095] = 32'hFFFFFFF1;
    // rom_array[14096] = 32'hFFFFFFF1;
    // rom_array[14097] = 32'hFFFFFFF0;
    // rom_array[14098] = 32'hFFFFFFF0;
    // rom_array[14099] = 32'hFFFFFFF0;
    // rom_array[14100] = 32'hFFFFFFF0;
    // rom_array[14101] = 32'hFFFFFFF1;
    // rom_array[14102] = 32'hFFFFFFF1;
    // rom_array[14103] = 32'hFFFFFFF1;
    // rom_array[14104] = 32'hFFFFFFF1;
    // rom_array[14105] = 32'hFFFFFFF0;
    // rom_array[14106] = 32'hFFFFFFF0;
    // rom_array[14107] = 32'hFFFFFFF0;
    // rom_array[14108] = 32'hFFFFFFF0;
    // rom_array[14109] = 32'hFFFFFFF1;
    // rom_array[14110] = 32'hFFFFFFF1;
    // rom_array[14111] = 32'hFFFFFFF1;
    // rom_array[14112] = 32'hFFFFFFF1;
    // rom_array[14113] = 32'hFFFFFFF0;
    // rom_array[14114] = 32'hFFFFFFF0;
    // rom_array[14115] = 32'hFFFFFFF0;
    // rom_array[14116] = 32'hFFFFFFF0;
    // rom_array[14117] = 32'hFFFFFFF1;
    // rom_array[14118] = 32'hFFFFFFF1;
    // rom_array[14119] = 32'hFFFFFFF1;
    // rom_array[14120] = 32'hFFFFFFF1;
    // rom_array[14121] = 32'hFFFFFFF0;
    // rom_array[14122] = 32'hFFFFFFF0;
    // rom_array[14123] = 32'hFFFFFFF0;
    // rom_array[14124] = 32'hFFFFFFF0;
    // rom_array[14125] = 32'hFFFFFFF1;
    // rom_array[14126] = 32'hFFFFFFF1;
    // rom_array[14127] = 32'hFFFFFFF1;
    // rom_array[14128] = 32'hFFFFFFF1;
    // rom_array[14129] = 32'hFFFFFFF0;
    // rom_array[14130] = 32'hFFFFFFF0;
    // rom_array[14131] = 32'hFFFFFFF0;
    // rom_array[14132] = 32'hFFFFFFF0;
    // rom_array[14133] = 32'hFFFFFFF1;
    // rom_array[14134] = 32'hFFFFFFF1;
    // rom_array[14135] = 32'hFFFFFFF1;
    // rom_array[14136] = 32'hFFFFFFF1;
    // rom_array[14137] = 32'hFFFFFFF0;
    // rom_array[14138] = 32'hFFFFFFF0;
    // rom_array[14139] = 32'hFFFFFFF0;
    // rom_array[14140] = 32'hFFFFFFF0;
    // rom_array[14141] = 32'hFFFFFFF1;
    // rom_array[14142] = 32'hFFFFFFF1;
    // rom_array[14143] = 32'hFFFFFFF1;
    // rom_array[14144] = 32'hFFFFFFF1;
    // rom_array[14145] = 32'hFFFFFFF0;
    // rom_array[14146] = 32'hFFFFFFF0;
    // rom_array[14147] = 32'hFFFFFFF0;
    // rom_array[14148] = 32'hFFFFFFF0;
    // rom_array[14149] = 32'hFFFFFFF1;
    // rom_array[14150] = 32'hFFFFFFF1;
    // rom_array[14151] = 32'hFFFFFFF1;
    // rom_array[14152] = 32'hFFFFFFF1;
    // rom_array[14153] = 32'hFFFFFFF0;
    // rom_array[14154] = 32'hFFFFFFF0;
    // rom_array[14155] = 32'hFFFFFFF0;
    // rom_array[14156] = 32'hFFFFFFF0;
    // rom_array[14157] = 32'hFFFFFFF1;
    // rom_array[14158] = 32'hFFFFFFF1;
    // rom_array[14159] = 32'hFFFFFFF1;
    // rom_array[14160] = 32'hFFFFFFF1;
    // rom_array[14161] = 32'hFFFFFFF0;
    // rom_array[14162] = 32'hFFFFFFF0;
    // rom_array[14163] = 32'hFFFFFFF0;
    // rom_array[14164] = 32'hFFFFFFF0;
    // rom_array[14165] = 32'hFFFFFFF1;
    // rom_array[14166] = 32'hFFFFFFF1;
    // rom_array[14167] = 32'hFFFFFFF1;
    // rom_array[14168] = 32'hFFFFFFF1;
    // rom_array[14169] = 32'hFFFFFFF0;
    // rom_array[14170] = 32'hFFFFFFF0;
    // rom_array[14171] = 32'hFFFFFFF0;
    // rom_array[14172] = 32'hFFFFFFF0;
    // rom_array[14173] = 32'hFFFFFFF1;
    // rom_array[14174] = 32'hFFFFFFF1;
    // rom_array[14175] = 32'hFFFFFFF1;
    // rom_array[14176] = 32'hFFFFFFF1;
    // rom_array[14177] = 32'hFFFFFFF0;
    // rom_array[14178] = 32'hFFFFFFF0;
    // rom_array[14179] = 32'hFFFFFFF0;
    // rom_array[14180] = 32'hFFFFFFF0;
    // rom_array[14181] = 32'hFFFFFFF1;
    // rom_array[14182] = 32'hFFFFFFF1;
    // rom_array[14183] = 32'hFFFFFFF1;
    // rom_array[14184] = 32'hFFFFFFF1;
    // rom_array[14185] = 32'hFFFFFFF1;
    // rom_array[14186] = 32'hFFFFFFF1;
    // rom_array[14187] = 32'hFFFFFFF1;
    // rom_array[14188] = 32'hFFFFFFF1;
    // rom_array[14189] = 32'hFFFFFFF1;
    // rom_array[14190] = 32'hFFFFFFF1;
    // rom_array[14191] = 32'hFFFFFFF1;
    // rom_array[14192] = 32'hFFFFFFF1;
    // rom_array[14193] = 32'hFFFFFFF1;
    // rom_array[14194] = 32'hFFFFFFF1;
    // rom_array[14195] = 32'hFFFFFFF1;
    // rom_array[14196] = 32'hFFFFFFF1;
    // rom_array[14197] = 32'hFFFFFFF1;
    // rom_array[14198] = 32'hFFFFFFF1;
    // rom_array[14199] = 32'hFFFFFFF1;
    // rom_array[14200] = 32'hFFFFFFF1;
    // rom_array[14201] = 32'hFFFFFFF0;
    // rom_array[14202] = 32'hFFFFFFF0;
    // rom_array[14203] = 32'hFFFFFFF0;
    // rom_array[14204] = 32'hFFFFFFF0;
    // rom_array[14205] = 32'hFFFFFFF1;
    // rom_array[14206] = 32'hFFFFFFF1;
    // rom_array[14207] = 32'hFFFFFFF1;
    // rom_array[14208] = 32'hFFFFFFF1;
    // rom_array[14209] = 32'hFFFFFFF0;
    // rom_array[14210] = 32'hFFFFFFF0;
    // rom_array[14211] = 32'hFFFFFFF0;
    // rom_array[14212] = 32'hFFFFFFF0;
    // rom_array[14213] = 32'hFFFFFFF1;
    // rom_array[14214] = 32'hFFFFFFF1;
    // rom_array[14215] = 32'hFFFFFFF1;
    // rom_array[14216] = 32'hFFFFFFF1;
    // rom_array[14217] = 32'hFFFFFFF0;
    // rom_array[14218] = 32'hFFFFFFF0;
    // rom_array[14219] = 32'hFFFFFFF0;
    // rom_array[14220] = 32'hFFFFFFF0;
    // rom_array[14221] = 32'hFFFFFFF1;
    // rom_array[14222] = 32'hFFFFFFF1;
    // rom_array[14223] = 32'hFFFFFFF1;
    // rom_array[14224] = 32'hFFFFFFF1;
    // rom_array[14225] = 32'hFFFFFFF0;
    // rom_array[14226] = 32'hFFFFFFF0;
    // rom_array[14227] = 32'hFFFFFFF0;
    // rom_array[14228] = 32'hFFFFFFF0;
    // rom_array[14229] = 32'hFFFFFFF1;
    // rom_array[14230] = 32'hFFFFFFF1;
    // rom_array[14231] = 32'hFFFFFFF1;
    // rom_array[14232] = 32'hFFFFFFF1;
    // rom_array[14233] = 32'hFFFFFFF1;
    // rom_array[14234] = 32'hFFFFFFF1;
    // rom_array[14235] = 32'hFFFFFFF1;
    // rom_array[14236] = 32'hFFFFFFF1;
    // rom_array[14237] = 32'hFFFFFFF1;
    // rom_array[14238] = 32'hFFFFFFF1;
    // rom_array[14239] = 32'hFFFFFFF1;
    // rom_array[14240] = 32'hFFFFFFF1;
    // rom_array[14241] = 32'hFFFFFFF1;
    // rom_array[14242] = 32'hFFFFFFF1;
    // rom_array[14243] = 32'hFFFFFFF1;
    // rom_array[14244] = 32'hFFFFFFF1;
    // rom_array[14245] = 32'hFFFFFFF1;
    // rom_array[14246] = 32'hFFFFFFF1;
    // rom_array[14247] = 32'hFFFFFFF1;
    // rom_array[14248] = 32'hFFFFFFF1;
    // rom_array[14249] = 32'hFFFFFFF1;
    // rom_array[14250] = 32'hFFFFFFF1;
    // rom_array[14251] = 32'hFFFFFFF1;
    // rom_array[14252] = 32'hFFFFFFF1;
    // rom_array[14253] = 32'hFFFFFFF1;
    // rom_array[14254] = 32'hFFFFFFF1;
    // rom_array[14255] = 32'hFFFFFFF1;
    // rom_array[14256] = 32'hFFFFFFF1;
    // rom_array[14257] = 32'hFFFFFFF1;
    // rom_array[14258] = 32'hFFFFFFF1;
    // rom_array[14259] = 32'hFFFFFFF1;
    // rom_array[14260] = 32'hFFFFFFF1;
    // rom_array[14261] = 32'hFFFFFFF1;
    // rom_array[14262] = 32'hFFFFFFF1;
    // rom_array[14263] = 32'hFFFFFFF1;
    // rom_array[14264] = 32'hFFFFFFF1;
    // rom_array[14265] = 32'hFFFFFFF0;
    // rom_array[14266] = 32'hFFFFFFF0;
    // rom_array[14267] = 32'hFFFFFFF0;
    // rom_array[14268] = 32'hFFFFFFF0;
    // rom_array[14269] = 32'hFFFFFFF1;
    // rom_array[14270] = 32'hFFFFFFF1;
    // rom_array[14271] = 32'hFFFFFFF1;
    // rom_array[14272] = 32'hFFFFFFF1;
    // rom_array[14273] = 32'hFFFFFFF0;
    // rom_array[14274] = 32'hFFFFFFF0;
    // rom_array[14275] = 32'hFFFFFFF0;
    // rom_array[14276] = 32'hFFFFFFF0;
    // rom_array[14277] = 32'hFFFFFFF1;
    // rom_array[14278] = 32'hFFFFFFF1;
    // rom_array[14279] = 32'hFFFFFFF1;
    // rom_array[14280] = 32'hFFFFFFF1;
    // rom_array[14281] = 32'hFFFFFFF0;
    // rom_array[14282] = 32'hFFFFFFF0;
    // rom_array[14283] = 32'hFFFFFFF0;
    // rom_array[14284] = 32'hFFFFFFF0;
    // rom_array[14285] = 32'hFFFFFFF1;
    // rom_array[14286] = 32'hFFFFFFF1;
    // rom_array[14287] = 32'hFFFFFFF1;
    // rom_array[14288] = 32'hFFFFFFF1;
    // rom_array[14289] = 32'hFFFFFFF0;
    // rom_array[14290] = 32'hFFFFFFF0;
    // rom_array[14291] = 32'hFFFFFFF0;
    // rom_array[14292] = 32'hFFFFFFF0;
    // rom_array[14293] = 32'hFFFFFFF1;
    // rom_array[14294] = 32'hFFFFFFF1;
    // rom_array[14295] = 32'hFFFFFFF1;
    // rom_array[14296] = 32'hFFFFFFF1;
    // rom_array[14297] = 32'hFFFFFFF1;
    // rom_array[14298] = 32'hFFFFFFF1;
    // rom_array[14299] = 32'hFFFFFFF1;
    // rom_array[14300] = 32'hFFFFFFF1;
    // rom_array[14301] = 32'hFFFFFFF1;
    // rom_array[14302] = 32'hFFFFFFF1;
    // rom_array[14303] = 32'hFFFFFFF1;
    // rom_array[14304] = 32'hFFFFFFF1;
    // rom_array[14305] = 32'hFFFFFFF1;
    // rom_array[14306] = 32'hFFFFFFF1;
    // rom_array[14307] = 32'hFFFFFFF1;
    // rom_array[14308] = 32'hFFFFFFF1;
    // rom_array[14309] = 32'hFFFFFFF1;
    // rom_array[14310] = 32'hFFFFFFF1;
    // rom_array[14311] = 32'hFFFFFFF1;
    // rom_array[14312] = 32'hFFFFFFF1;
    // rom_array[14313] = 32'hFFFFFFF1;
    // rom_array[14314] = 32'hFFFFFFF1;
    // rom_array[14315] = 32'hFFFFFFF1;
    // rom_array[14316] = 32'hFFFFFFF1;
    // rom_array[14317] = 32'hFFFFFFF1;
    // rom_array[14318] = 32'hFFFFFFF1;
    // rom_array[14319] = 32'hFFFFFFF1;
    // rom_array[14320] = 32'hFFFFFFF1;
    // rom_array[14321] = 32'hFFFFFFF1;
    // rom_array[14322] = 32'hFFFFFFF1;
    // rom_array[14323] = 32'hFFFFFFF1;
    // rom_array[14324] = 32'hFFFFFFF1;
    // rom_array[14325] = 32'hFFFFFFF1;
    // rom_array[14326] = 32'hFFFFFFF1;
    // rom_array[14327] = 32'hFFFFFFF1;
    // rom_array[14328] = 32'hFFFFFFF1;
    // rom_array[14329] = 32'hFFFFFFF0;
    // rom_array[14330] = 32'hFFFFFFF0;
    // rom_array[14331] = 32'hFFFFFFF1;
    // rom_array[14332] = 32'hFFFFFFF1;
    // rom_array[14333] = 32'hFFFFFFF0;
    // rom_array[14334] = 32'hFFFFFFF0;
    // rom_array[14335] = 32'hFFFFFFF1;
    // rom_array[14336] = 32'hFFFFFFF1;
    // rom_array[14337] = 32'hFFFFFFF0;
    // rom_array[14338] = 32'hFFFFFFF0;
    // rom_array[14339] = 32'hFFFFFFF1;
    // rom_array[14340] = 32'hFFFFFFF1;
    // rom_array[14341] = 32'hFFFFFFF0;
    // rom_array[14342] = 32'hFFFFFFF0;
    // rom_array[14343] = 32'hFFFFFFF1;
    // rom_array[14344] = 32'hFFFFFFF1;
    // rom_array[14345] = 32'hFFFFFFF0;
    // rom_array[14346] = 32'hFFFFFFF0;
    // rom_array[14347] = 32'hFFFFFFF1;
    // rom_array[14348] = 32'hFFFFFFF1;
    // rom_array[14349] = 32'hFFFFFFF0;
    // rom_array[14350] = 32'hFFFFFFF0;
    // rom_array[14351] = 32'hFFFFFFF1;
    // rom_array[14352] = 32'hFFFFFFF1;
    // rom_array[14353] = 32'hFFFFFFF0;
    // rom_array[14354] = 32'hFFFFFFF0;
    // rom_array[14355] = 32'hFFFFFFF1;
    // rom_array[14356] = 32'hFFFFFFF1;
    // rom_array[14357] = 32'hFFFFFFF0;
    // rom_array[14358] = 32'hFFFFFFF0;
    // rom_array[14359] = 32'hFFFFFFF1;
    // rom_array[14360] = 32'hFFFFFFF1;
    // rom_array[14361] = 32'hFFFFFFF0;
    // rom_array[14362] = 32'hFFFFFFF0;
    // rom_array[14363] = 32'hFFFFFFF1;
    // rom_array[14364] = 32'hFFFFFFF1;
    // rom_array[14365] = 32'hFFFFFFF0;
    // rom_array[14366] = 32'hFFFFFFF0;
    // rom_array[14367] = 32'hFFFFFFF0;
    // rom_array[14368] = 32'hFFFFFFF0;
    // rom_array[14369] = 32'hFFFFFFF0;
    // rom_array[14370] = 32'hFFFFFFF0;
    // rom_array[14371] = 32'hFFFFFFF1;
    // rom_array[14372] = 32'hFFFFFFF1;
    // rom_array[14373] = 32'hFFFFFFF0;
    // rom_array[14374] = 32'hFFFFFFF0;
    // rom_array[14375] = 32'hFFFFFFF0;
    // rom_array[14376] = 32'hFFFFFFF0;
    // rom_array[14377] = 32'hFFFFFFF1;
    // rom_array[14378] = 32'hFFFFFFF1;
    // rom_array[14379] = 32'hFFFFFFF1;
    // rom_array[14380] = 32'hFFFFFFF1;
    // rom_array[14381] = 32'hFFFFFFF0;
    // rom_array[14382] = 32'hFFFFFFF0;
    // rom_array[14383] = 32'hFFFFFFF0;
    // rom_array[14384] = 32'hFFFFFFF0;
    // rom_array[14385] = 32'hFFFFFFF1;
    // rom_array[14386] = 32'hFFFFFFF1;
    // rom_array[14387] = 32'hFFFFFFF1;
    // rom_array[14388] = 32'hFFFFFFF1;
    // rom_array[14389] = 32'hFFFFFFF0;
    // rom_array[14390] = 32'hFFFFFFF0;
    // rom_array[14391] = 32'hFFFFFFF0;
    // rom_array[14392] = 32'hFFFFFFF0;
    // rom_array[14393] = 32'hFFFFFFF1;
    // rom_array[14394] = 32'hFFFFFFF1;
    // rom_array[14395] = 32'hFFFFFFF1;
    // rom_array[14396] = 32'hFFFFFFF1;
    // rom_array[14397] = 32'hFFFFFFF0;
    // rom_array[14398] = 32'hFFFFFFF0;
    // rom_array[14399] = 32'hFFFFFFF0;
    // rom_array[14400] = 32'hFFFFFFF0;
    // rom_array[14401] = 32'hFFFFFFF1;
    // rom_array[14402] = 32'hFFFFFFF1;
    // rom_array[14403] = 32'hFFFFFFF1;
    // rom_array[14404] = 32'hFFFFFFF1;
    // rom_array[14405] = 32'hFFFFFFF0;
    // rom_array[14406] = 32'hFFFFFFF0;
    // rom_array[14407] = 32'hFFFFFFF0;
    // rom_array[14408] = 32'hFFFFFFF0;
    // rom_array[14409] = 32'hFFFFFFF1;
    // rom_array[14410] = 32'hFFFFFFF1;
    // rom_array[14411] = 32'hFFFFFFF1;
    // rom_array[14412] = 32'hFFFFFFF1;
    // rom_array[14413] = 32'hFFFFFFF0;
    // rom_array[14414] = 32'hFFFFFFF0;
    // rom_array[14415] = 32'hFFFFFFF0;
    // rom_array[14416] = 32'hFFFFFFF0;
    // rom_array[14417] = 32'hFFFFFFF1;
    // rom_array[14418] = 32'hFFFFFFF1;
    // rom_array[14419] = 32'hFFFFFFF1;
    // rom_array[14420] = 32'hFFFFFFF1;
    // rom_array[14421] = 32'hFFFFFFF0;
    // rom_array[14422] = 32'hFFFFFFF0;
    // rom_array[14423] = 32'hFFFFFFF0;
    // rom_array[14424] = 32'hFFFFFFF0;
    // rom_array[14425] = 32'hFFFFFFF1;
    // rom_array[14426] = 32'hFFFFFFF1;
    // rom_array[14427] = 32'hFFFFFFF1;
    // rom_array[14428] = 32'hFFFFFFF1;
    // rom_array[14429] = 32'hFFFFFFF1;
    // rom_array[14430] = 32'hFFFFFFF1;
    // rom_array[14431] = 32'hFFFFFFF1;
    // rom_array[14432] = 32'hFFFFFFF1;
    // rom_array[14433] = 32'hFFFFFFF1;
    // rom_array[14434] = 32'hFFFFFFF1;
    // rom_array[14435] = 32'hFFFFFFF1;
    // rom_array[14436] = 32'hFFFFFFF1;
    // rom_array[14437] = 32'hFFFFFFF1;
    // rom_array[14438] = 32'hFFFFFFF1;
    // rom_array[14439] = 32'hFFFFFFF1;
    // rom_array[14440] = 32'hFFFFFFF1;
    // rom_array[14441] = 32'hFFFFFFF1;
    // rom_array[14442] = 32'hFFFFFFF1;
    // rom_array[14443] = 32'hFFFFFFF1;
    // rom_array[14444] = 32'hFFFFFFF1;
    // rom_array[14445] = 32'hFFFFFFF1;
    // rom_array[14446] = 32'hFFFFFFF1;
    // rom_array[14447] = 32'hFFFFFFF1;
    // rom_array[14448] = 32'hFFFFFFF1;
    // rom_array[14449] = 32'hFFFFFFF1;
    // rom_array[14450] = 32'hFFFFFFF1;
    // rom_array[14451] = 32'hFFFFFFF1;
    // rom_array[14452] = 32'hFFFFFFF1;
    // rom_array[14453] = 32'hFFFFFFF1;
    // rom_array[14454] = 32'hFFFFFFF1;
    // rom_array[14455] = 32'hFFFFFFF1;
    // rom_array[14456] = 32'hFFFFFFF1;
    // rom_array[14457] = 32'hFFFFFFF1;
    // rom_array[14458] = 32'hFFFFFFF1;
    // rom_array[14459] = 32'hFFFFFFF1;
    // rom_array[14460] = 32'hFFFFFFF1;
    // rom_array[14461] = 32'hFFFFFFF0;
    // rom_array[14462] = 32'hFFFFFFF0;
    // rom_array[14463] = 32'hFFFFFFF0;
    // rom_array[14464] = 32'hFFFFFFF0;
    // rom_array[14465] = 32'hFFFFFFF1;
    // rom_array[14466] = 32'hFFFFFFF1;
    // rom_array[14467] = 32'hFFFFFFF1;
    // rom_array[14468] = 32'hFFFFFFF1;
    // rom_array[14469] = 32'hFFFFFFF0;
    // rom_array[14470] = 32'hFFFFFFF0;
    // rom_array[14471] = 32'hFFFFFFF0;
    // rom_array[14472] = 32'hFFFFFFF0;
    // rom_array[14473] = 32'hFFFFFFF1;
    // rom_array[14474] = 32'hFFFFFFF1;
    // rom_array[14475] = 32'hFFFFFFF1;
    // rom_array[14476] = 32'hFFFFFFF1;
    // rom_array[14477] = 32'hFFFFFFF0;
    // rom_array[14478] = 32'hFFFFFFF0;
    // rom_array[14479] = 32'hFFFFFFF0;
    // rom_array[14480] = 32'hFFFFFFF0;
    // rom_array[14481] = 32'hFFFFFFF1;
    // rom_array[14482] = 32'hFFFFFFF1;
    // rom_array[14483] = 32'hFFFFFFF1;
    // rom_array[14484] = 32'hFFFFFFF1;
    // rom_array[14485] = 32'hFFFFFFF0;
    // rom_array[14486] = 32'hFFFFFFF0;
    // rom_array[14487] = 32'hFFFFFFF0;
    // rom_array[14488] = 32'hFFFFFFF0;
    // rom_array[14489] = 32'hFFFFFFF1;
    // rom_array[14490] = 32'hFFFFFFF1;
    // rom_array[14491] = 32'hFFFFFFF1;
    // rom_array[14492] = 32'hFFFFFFF1;
    // rom_array[14493] = 32'hFFFFFFF0;
    // rom_array[14494] = 32'hFFFFFFF0;
    // rom_array[14495] = 32'hFFFFFFF0;
    // rom_array[14496] = 32'hFFFFFFF0;
    // rom_array[14497] = 32'hFFFFFFF1;
    // rom_array[14498] = 32'hFFFFFFF1;
    // rom_array[14499] = 32'hFFFFFFF1;
    // rom_array[14500] = 32'hFFFFFFF1;
    // rom_array[14501] = 32'hFFFFFFF0;
    // rom_array[14502] = 32'hFFFFFFF0;
    // rom_array[14503] = 32'hFFFFFFF0;
    // rom_array[14504] = 32'hFFFFFFF0;
    // rom_array[14505] = 32'hFFFFFFF1;
    // rom_array[14506] = 32'hFFFFFFF1;
    // rom_array[14507] = 32'hFFFFFFF1;
    // rom_array[14508] = 32'hFFFFFFF1;
    // rom_array[14509] = 32'hFFFFFFF1;
    // rom_array[14510] = 32'hFFFFFFF1;
    // rom_array[14511] = 32'hFFFFFFF1;
    // rom_array[14512] = 32'hFFFFFFF1;
    // rom_array[14513] = 32'hFFFFFFF1;
    // rom_array[14514] = 32'hFFFFFFF1;
    // rom_array[14515] = 32'hFFFFFFF1;
    // rom_array[14516] = 32'hFFFFFFF1;
    // rom_array[14517] = 32'hFFFFFFF1;
    // rom_array[14518] = 32'hFFFFFFF1;
    // rom_array[14519] = 32'hFFFFFFF1;
    // rom_array[14520] = 32'hFFFFFFF1;
    // rom_array[14521] = 32'hFFFFFFF1;
    // rom_array[14522] = 32'hFFFFFFF1;
    // rom_array[14523] = 32'hFFFFFFF1;
    // rom_array[14524] = 32'hFFFFFFF1;
    // rom_array[14525] = 32'hFFFFFFF1;
    // rom_array[14526] = 32'hFFFFFFF1;
    // rom_array[14527] = 32'hFFFFFFF1;
    // rom_array[14528] = 32'hFFFFFFF1;
    // rom_array[14529] = 32'hFFFFFFF1;
    // rom_array[14530] = 32'hFFFFFFF1;
    // rom_array[14531] = 32'hFFFFFFF1;
    // rom_array[14532] = 32'hFFFFFFF1;
    // rom_array[14533] = 32'hFFFFFFF1;
    // rom_array[14534] = 32'hFFFFFFF1;
    // rom_array[14535] = 32'hFFFFFFF1;
    // rom_array[14536] = 32'hFFFFFFF1;
    // rom_array[14537] = 32'hFFFFFFF1;
    // rom_array[14538] = 32'hFFFFFFF1;
    // rom_array[14539] = 32'hFFFFFFF1;
    // rom_array[14540] = 32'hFFFFFFF1;
    // rom_array[14541] = 32'hFFFFFFF0;
    // rom_array[14542] = 32'hFFFFFFF0;
    // rom_array[14543] = 32'hFFFFFFF0;
    // rom_array[14544] = 32'hFFFFFFF0;
    // rom_array[14545] = 32'hFFFFFFF1;
    // rom_array[14546] = 32'hFFFFFFF1;
    // rom_array[14547] = 32'hFFFFFFF1;
    // rom_array[14548] = 32'hFFFFFFF1;
    // rom_array[14549] = 32'hFFFFFFF0;
    // rom_array[14550] = 32'hFFFFFFF0;
    // rom_array[14551] = 32'hFFFFFFF0;
    // rom_array[14552] = 32'hFFFFFFF0;
    // rom_array[14553] = 32'hFFFFFFF1;
    // rom_array[14554] = 32'hFFFFFFF1;
    // rom_array[14555] = 32'hFFFFFFF1;
    // rom_array[14556] = 32'hFFFFFFF1;
    // rom_array[14557] = 32'hFFFFFFF0;
    // rom_array[14558] = 32'hFFFFFFF0;
    // rom_array[14559] = 32'hFFFFFFF0;
    // rom_array[14560] = 32'hFFFFFFF0;
    // rom_array[14561] = 32'hFFFFFFF1;
    // rom_array[14562] = 32'hFFFFFFF1;
    // rom_array[14563] = 32'hFFFFFFF1;
    // rom_array[14564] = 32'hFFFFFFF1;
    // rom_array[14565] = 32'hFFFFFFF0;
    // rom_array[14566] = 32'hFFFFFFF0;
    // rom_array[14567] = 32'hFFFFFFF0;
    // rom_array[14568] = 32'hFFFFFFF0;
    // rom_array[14569] = 32'hFFFFFFF1;
    // rom_array[14570] = 32'hFFFFFFF1;
    // rom_array[14571] = 32'hFFFFFFF1;
    // rom_array[14572] = 32'hFFFFFFF1;
    // rom_array[14573] = 32'hFFFFFFF0;
    // rom_array[14574] = 32'hFFFFFFF0;
    // rom_array[14575] = 32'hFFFFFFF0;
    // rom_array[14576] = 32'hFFFFFFF0;
    // rom_array[14577] = 32'hFFFFFFF1;
    // rom_array[14578] = 32'hFFFFFFF1;
    // rom_array[14579] = 32'hFFFFFFF1;
    // rom_array[14580] = 32'hFFFFFFF1;
    // rom_array[14581] = 32'hFFFFFFF0;
    // rom_array[14582] = 32'hFFFFFFF0;
    // rom_array[14583] = 32'hFFFFFFF0;
    // rom_array[14584] = 32'hFFFFFFF0;
    // rom_array[14585] = 32'hFFFFFFF1;
    // rom_array[14586] = 32'hFFFFFFF1;
    // rom_array[14587] = 32'hFFFFFFF1;
    // rom_array[14588] = 32'hFFFFFFF1;
    // rom_array[14589] = 32'hFFFFFFF0;
    // rom_array[14590] = 32'hFFFFFFF0;
    // rom_array[14591] = 32'hFFFFFFF0;
    // rom_array[14592] = 32'hFFFFFFF0;
    // rom_array[14593] = 32'hFFFFFFF1;
    // rom_array[14594] = 32'hFFFFFFF1;
    // rom_array[14595] = 32'hFFFFFFF1;
    // rom_array[14596] = 32'hFFFFFFF1;
    // rom_array[14597] = 32'hFFFFFFF0;
    // rom_array[14598] = 32'hFFFFFFF0;
    // rom_array[14599] = 32'hFFFFFFF0;
    // rom_array[14600] = 32'hFFFFFFF0;
    // rom_array[14601] = 32'hFFFFFFF1;
    // rom_array[14602] = 32'hFFFFFFF1;
    // rom_array[14603] = 32'hFFFFFFF1;
    // rom_array[14604] = 32'hFFFFFFF1;
    // rom_array[14605] = 32'hFFFFFFF1;
    // rom_array[14606] = 32'hFFFFFFF1;
    // rom_array[14607] = 32'hFFFFFFF1;
    // rom_array[14608] = 32'hFFFFFFF1;
    // rom_array[14609] = 32'hFFFFFFF1;
    // rom_array[14610] = 32'hFFFFFFF1;
    // rom_array[14611] = 32'hFFFFFFF1;
    // rom_array[14612] = 32'hFFFFFFF1;
    // rom_array[14613] = 32'hFFFFFFF1;
    // rom_array[14614] = 32'hFFFFFFF1;
    // rom_array[14615] = 32'hFFFFFFF1;
    // rom_array[14616] = 32'hFFFFFFF1;
    // rom_array[14617] = 32'hFFFFFFF1;
    // rom_array[14618] = 32'hFFFFFFF1;
    // rom_array[14619] = 32'hFFFFFFF1;
    // rom_array[14620] = 32'hFFFFFFF1;
    // rom_array[14621] = 32'hFFFFFFF1;
    // rom_array[14622] = 32'hFFFFFFF1;
    // rom_array[14623] = 32'hFFFFFFF1;
    // rom_array[14624] = 32'hFFFFFFF1;
    // rom_array[14625] = 32'hFFFFFFF1;
    // rom_array[14626] = 32'hFFFFFFF1;
    // rom_array[14627] = 32'hFFFFFFF1;
    // rom_array[14628] = 32'hFFFFFFF1;
    // rom_array[14629] = 32'hFFFFFFF1;
    // rom_array[14630] = 32'hFFFFFFF1;
    // rom_array[14631] = 32'hFFFFFFF1;
    // rom_array[14632] = 32'hFFFFFFF1;
    // rom_array[14633] = 32'hFFFFFFF1;
    // rom_array[14634] = 32'hFFFFFFF1;
    // rom_array[14635] = 32'hFFFFFFF1;
    // rom_array[14636] = 32'hFFFFFFF1;
    // rom_array[14637] = 32'hFFFFFFF1;
    // rom_array[14638] = 32'hFFFFFFF1;
    // rom_array[14639] = 32'hFFFFFFF1;
    // rom_array[14640] = 32'hFFFFFFF1;
    // rom_array[14641] = 32'hFFFFFFF1;
    // rom_array[14642] = 32'hFFFFFFF1;
    // rom_array[14643] = 32'hFFFFFFF1;
    // rom_array[14644] = 32'hFFFFFFF1;
    // rom_array[14645] = 32'hFFFFFFF1;
    // rom_array[14646] = 32'hFFFFFFF1;
    // rom_array[14647] = 32'hFFFFFFF1;
    // rom_array[14648] = 32'hFFFFFFF1;
    // rom_array[14649] = 32'hFFFFFFF1;
    // rom_array[14650] = 32'hFFFFFFF1;
    // rom_array[14651] = 32'hFFFFFFF1;
    // rom_array[14652] = 32'hFFFFFFF1;
    // rom_array[14653] = 32'hFFFFFFF1;
    // rom_array[14654] = 32'hFFFFFFF1;
    // rom_array[14655] = 32'hFFFFFFF1;
    // rom_array[14656] = 32'hFFFFFFF1;
    // rom_array[14657] = 32'hFFFFFFF1;
    // rom_array[14658] = 32'hFFFFFFF1;
    // rom_array[14659] = 32'hFFFFFFF1;
    // rom_array[14660] = 32'hFFFFFFF1;
    // rom_array[14661] = 32'hFFFFFFF1;
    // rom_array[14662] = 32'hFFFFFFF1;
    // rom_array[14663] = 32'hFFFFFFF1;
    // rom_array[14664] = 32'hFFFFFFF1;
    // rom_array[14665] = 32'hFFFFFFF1;
    // rom_array[14666] = 32'hFFFFFFF1;
    // rom_array[14667] = 32'hFFFFFFF1;
    // rom_array[14668] = 32'hFFFFFFF1;
    // rom_array[14669] = 32'hFFFFFFF1;
    // rom_array[14670] = 32'hFFFFFFF1;
    // rom_array[14671] = 32'hFFFFFFF1;
    // rom_array[14672] = 32'hFFFFFFF1;
    // rom_array[14673] = 32'hFFFFFFF1;
    // rom_array[14674] = 32'hFFFFFFF1;
    // rom_array[14675] = 32'hFFFFFFF1;
    // rom_array[14676] = 32'hFFFFFFF1;
    // rom_array[14677] = 32'hFFFFFFF1;
    // rom_array[14678] = 32'hFFFFFFF1;
    // rom_array[14679] = 32'hFFFFFFF1;
    // rom_array[14680] = 32'hFFFFFFF1;
    // rom_array[14681] = 32'hFFFFFFF1;
    // rom_array[14682] = 32'hFFFFFFF1;
    // rom_array[14683] = 32'hFFFFFFF1;
    // rom_array[14684] = 32'hFFFFFFF1;
    // rom_array[14685] = 32'hFFFFFFF1;
    // rom_array[14686] = 32'hFFFFFFF1;
    // rom_array[14687] = 32'hFFFFFFF1;
    // rom_array[14688] = 32'hFFFFFFF1;
    // rom_array[14689] = 32'hFFFFFFF1;
    // rom_array[14690] = 32'hFFFFFFF1;
    // rom_array[14691] = 32'hFFFFFFF1;
    // rom_array[14692] = 32'hFFFFFFF1;
    // rom_array[14693] = 32'hFFFFFFF1;
    // rom_array[14694] = 32'hFFFFFFF1;
    // rom_array[14695] = 32'hFFFFFFF1;
    // rom_array[14696] = 32'hFFFFFFF1;
    // rom_array[14697] = 32'hFFFFFFF1;
    // rom_array[14698] = 32'hFFFFFFF1;
    // rom_array[14699] = 32'hFFFFFFF1;
    // rom_array[14700] = 32'hFFFFFFF1;
    // rom_array[14701] = 32'hFFFFFFF1;
    // rom_array[14702] = 32'hFFFFFFF1;
    // rom_array[14703] = 32'hFFFFFFF1;
    // rom_array[14704] = 32'hFFFFFFF1;
    // rom_array[14705] = 32'hFFFFFFF1;
    // rom_array[14706] = 32'hFFFFFFF1;
    // rom_array[14707] = 32'hFFFFFFF1;
    // rom_array[14708] = 32'hFFFFFFF1;
    // rom_array[14709] = 32'hFFFFFFF1;
    // rom_array[14710] = 32'hFFFFFFF1;
    // rom_array[14711] = 32'hFFFFFFF1;
    // rom_array[14712] = 32'hFFFFFFF1;
    // rom_array[14713] = 32'hFFFFFFF1;
    // rom_array[14714] = 32'hFFFFFFF1;
    // rom_array[14715] = 32'hFFFFFFF1;
    // rom_array[14716] = 32'hFFFFFFF1;
    // rom_array[14717] = 32'hFFFFFFF1;
    // rom_array[14718] = 32'hFFFFFFF1;
    // rom_array[14719] = 32'hFFFFFFF1;
    // rom_array[14720] = 32'hFFFFFFF1;
    // rom_array[14721] = 32'hFFFFFFF1;
    // rom_array[14722] = 32'hFFFFFFF1;
    // rom_array[14723] = 32'hFFFFFFF1;
    // rom_array[14724] = 32'hFFFFFFF1;
    // rom_array[14725] = 32'hFFFFFFF1;
    // rom_array[14726] = 32'hFFFFFFF1;
    // rom_array[14727] = 32'hFFFFFFF1;
    // rom_array[14728] = 32'hFFFFFFF1;
    // rom_array[14729] = 32'hFFFFFFF1;
    // rom_array[14730] = 32'hFFFFFFF1;
    // rom_array[14731] = 32'hFFFFFFF1;
    // rom_array[14732] = 32'hFFFFFFF1;
    // rom_array[14733] = 32'hFFFFFFF1;
    // rom_array[14734] = 32'hFFFFFFF1;
    // rom_array[14735] = 32'hFFFFFFF1;
    // rom_array[14736] = 32'hFFFFFFF1;
    // rom_array[14737] = 32'hFFFFFFF1;
    // rom_array[14738] = 32'hFFFFFFF1;
    // rom_array[14739] = 32'hFFFFFFF1;
    // rom_array[14740] = 32'hFFFFFFF1;
    // rom_array[14741] = 32'hFFFFFFF1;
    // rom_array[14742] = 32'hFFFFFFF1;
    // rom_array[14743] = 32'hFFFFFFF1;
    // rom_array[14744] = 32'hFFFFFFF1;
    // rom_array[14745] = 32'hFFFFFFF1;
    // rom_array[14746] = 32'hFFFFFFF1;
    // rom_array[14747] = 32'hFFFFFFF1;
    // rom_array[14748] = 32'hFFFFFFF1;
    // rom_array[14749] = 32'hFFFFFFF1;
    // rom_array[14750] = 32'hFFFFFFF1;
    // rom_array[14751] = 32'hFFFFFFF1;
    // rom_array[14752] = 32'hFFFFFFF1;
    // rom_array[14753] = 32'hFFFFFFF1;
    // rom_array[14754] = 32'hFFFFFFF1;
    // rom_array[14755] = 32'hFFFFFFF1;
    // rom_array[14756] = 32'hFFFFFFF1;
    // rom_array[14757] = 32'hFFFFFFF1;
    // rom_array[14758] = 32'hFFFFFFF1;
    // rom_array[14759] = 32'hFFFFFFF1;
    // rom_array[14760] = 32'hFFFFFFF1;
    // rom_array[14761] = 32'hFFFFFFF1;
    // rom_array[14762] = 32'hFFFFFFF1;
    // rom_array[14763] = 32'hFFFFFFF1;
    // rom_array[14764] = 32'hFFFFFFF1;
    // rom_array[14765] = 32'hFFFFFFF1;
    // rom_array[14766] = 32'hFFFFFFF1;
    // rom_array[14767] = 32'hFFFFFFF1;
    // rom_array[14768] = 32'hFFFFFFF1;
    // rom_array[14769] = 32'hFFFFFFF1;
    // rom_array[14770] = 32'hFFFFFFF1;
    // rom_array[14771] = 32'hFFFFFFF1;
    // rom_array[14772] = 32'hFFFFFFF1;
    // rom_array[14773] = 32'hFFFFFFF1;
    // rom_array[14774] = 32'hFFFFFFF1;
    // rom_array[14775] = 32'hFFFFFFF1;
    // rom_array[14776] = 32'hFFFFFFF1;
    // rom_array[14777] = 32'hFFFFFFF1;
    // rom_array[14778] = 32'hFFFFFFF1;
    // rom_array[14779] = 32'hFFFFFFF1;
    // rom_array[14780] = 32'hFFFFFFF1;
    // rom_array[14781] = 32'hFFFFFFF1;
    // rom_array[14782] = 32'hFFFFFFF1;
    // rom_array[14783] = 32'hFFFFFFF1;
    // rom_array[14784] = 32'hFFFFFFF1;
    // rom_array[14785] = 32'hFFFFFFF1;
    // rom_array[14786] = 32'hFFFFFFF1;
    // rom_array[14787] = 32'hFFFFFFF1;
    // rom_array[14788] = 32'hFFFFFFF1;
    // rom_array[14789] = 32'hFFFFFFF1;
    // rom_array[14790] = 32'hFFFFFFF1;
    // rom_array[14791] = 32'hFFFFFFF1;
    // rom_array[14792] = 32'hFFFFFFF1;
    // rom_array[14793] = 32'hFFFFFFF1;
    // rom_array[14794] = 32'hFFFFFFF1;
    // rom_array[14795] = 32'hFFFFFFF1;
    // rom_array[14796] = 32'hFFFFFFF1;
    // rom_array[14797] = 32'hFFFFFFF1;
    // rom_array[14798] = 32'hFFFFFFF1;
    // rom_array[14799] = 32'hFFFFFFF1;
    // rom_array[14800] = 32'hFFFFFFF1;
    // rom_array[14801] = 32'hFFFFFFF1;
    // rom_array[14802] = 32'hFFFFFFF1;
    // rom_array[14803] = 32'hFFFFFFF1;
    // rom_array[14804] = 32'hFFFFFFF1;
    // rom_array[14805] = 32'hFFFFFFF1;
    // rom_array[14806] = 32'hFFFFFFF1;
    // rom_array[14807] = 32'hFFFFFFF1;
    // rom_array[14808] = 32'hFFFFFFF1;
    // rom_array[14809] = 32'hFFFFFFF1;
    // rom_array[14810] = 32'hFFFFFFF1;
    // rom_array[14811] = 32'hFFFFFFF1;
    // rom_array[14812] = 32'hFFFFFFF1;
    // rom_array[14813] = 32'hFFFFFFF1;
    // rom_array[14814] = 32'hFFFFFFF1;
    // rom_array[14815] = 32'hFFFFFFF1;
    // rom_array[14816] = 32'hFFFFFFF1;
    // rom_array[14817] = 32'hFFFFFFF1;
    // rom_array[14818] = 32'hFFFFFFF1;
    // rom_array[14819] = 32'hFFFFFFF1;
    // rom_array[14820] = 32'hFFFFFFF1;
    // rom_array[14821] = 32'hFFFFFFF1;
    // rom_array[14822] = 32'hFFFFFFF1;
    // rom_array[14823] = 32'hFFFFFFF1;
    // rom_array[14824] = 32'hFFFFFFF1;
    // rom_array[14825] = 32'hFFFFFFF1;
    // rom_array[14826] = 32'hFFFFFFF1;
    // rom_array[14827] = 32'hFFFFFFF1;
    // rom_array[14828] = 32'hFFFFFFF1;
    // rom_array[14829] = 32'hFFFFFFF1;
    // rom_array[14830] = 32'hFFFFFFF1;
    // rom_array[14831] = 32'hFFFFFFF1;
    // rom_array[14832] = 32'hFFFFFFF1;
    // rom_array[14833] = 32'hFFFFFFF1;
    // rom_array[14834] = 32'hFFFFFFF1;
    // rom_array[14835] = 32'hFFFFFFF1;
    // rom_array[14836] = 32'hFFFFFFF1;
    // rom_array[14837] = 32'hFFFFFFF1;
    // rom_array[14838] = 32'hFFFFFFF1;
    // rom_array[14839] = 32'hFFFFFFF1;
    // rom_array[14840] = 32'hFFFFFFF1;
    // rom_array[14841] = 32'hFFFFFFF1;
    // rom_array[14842] = 32'hFFFFFFF1;
    // rom_array[14843] = 32'hFFFFFFF1;
    // rom_array[14844] = 32'hFFFFFFF1;
    // rom_array[14845] = 32'hFFFFFFF1;
    // rom_array[14846] = 32'hFFFFFFF1;
    // rom_array[14847] = 32'hFFFFFFF1;
    // rom_array[14848] = 32'hFFFFFFF1;
    // rom_array[14849] = 32'hFFFFFFF1;
    // rom_array[14850] = 32'hFFFFFFF1;
    // rom_array[14851] = 32'hFFFFFFF1;
    // rom_array[14852] = 32'hFFFFFFF1;
    // rom_array[14853] = 32'hFFFFFFF1;
    // rom_array[14854] = 32'hFFFFFFF1;
    // rom_array[14855] = 32'hFFFFFFF1;
    // rom_array[14856] = 32'hFFFFFFF1;
    // rom_array[14857] = 32'hFFFFFFF1;
    // rom_array[14858] = 32'hFFFFFFF1;
    // rom_array[14859] = 32'hFFFFFFF1;
    // rom_array[14860] = 32'hFFFFFFF1;
    // rom_array[14861] = 32'hFFFFFFF1;
    // rom_array[14862] = 32'hFFFFFFF1;
    // rom_array[14863] = 32'hFFFFFFF1;
    // rom_array[14864] = 32'hFFFFFFF1;
    // rom_array[14865] = 32'hFFFFFFF1;
    // rom_array[14866] = 32'hFFFFFFF1;
    // rom_array[14867] = 32'hFFFFFFF1;
    // rom_array[14868] = 32'hFFFFFFF1;
    // rom_array[14869] = 32'hFFFFFFF1;
    // rom_array[14870] = 32'hFFFFFFF1;
    // rom_array[14871] = 32'hFFFFFFF1;
    // rom_array[14872] = 32'hFFFFFFF1;
    // rom_array[14873] = 32'hFFFFFFF1;
    // rom_array[14874] = 32'hFFFFFFF1;
    // rom_array[14875] = 32'hFFFFFFF1;
    // rom_array[14876] = 32'hFFFFFFF1;
    // rom_array[14877] = 32'hFFFFFFF1;
    // rom_array[14878] = 32'hFFFFFFF1;
    // rom_array[14879] = 32'hFFFFFFF1;
    // rom_array[14880] = 32'hFFFFFFF1;
    // rom_array[14881] = 32'hFFFFFFF1;
    // rom_array[14882] = 32'hFFFFFFF1;
    // rom_array[14883] = 32'hFFFFFFF1;
    // rom_array[14884] = 32'hFFFFFFF1;
    // rom_array[14885] = 32'hFFFFFFF1;
    // rom_array[14886] = 32'hFFFFFFF1;
    // rom_array[14887] = 32'hFFFFFFF1;
    // rom_array[14888] = 32'hFFFFFFF1;
    // rom_array[14889] = 32'hFFFFFFF1;
    // rom_array[14890] = 32'hFFFFFFF1;
    // rom_array[14891] = 32'hFFFFFFF1;
    // rom_array[14892] = 32'hFFFFFFF1;
    // rom_array[14893] = 32'hFFFFFFF1;
    // rom_array[14894] = 32'hFFFFFFF1;
    // rom_array[14895] = 32'hFFFFFFF1;
    // rom_array[14896] = 32'hFFFFFFF1;
    // rom_array[14897] = 32'hFFFFFFF1;
    // rom_array[14898] = 32'hFFFFFFF1;
    // rom_array[14899] = 32'hFFFFFFF1;
    // rom_array[14900] = 32'hFFFFFFF1;
    // rom_array[14901] = 32'hFFFFFFF1;
    // rom_array[14902] = 32'hFFFFFFF1;
    // rom_array[14903] = 32'hFFFFFFF1;
    // rom_array[14904] = 32'hFFFFFFF1;
    // rom_array[14905] = 32'hFFFFFFF1;
    // rom_array[14906] = 32'hFFFFFFF1;
    // rom_array[14907] = 32'hFFFFFFF1;
    // rom_array[14908] = 32'hFFFFFFF1;
    // rom_array[14909] = 32'hFFFFFFF1;
    // rom_array[14910] = 32'hFFFFFFF1;
    // rom_array[14911] = 32'hFFFFFFF1;
    // rom_array[14912] = 32'hFFFFFFF1;
    // rom_array[14913] = 32'hFFFFFFF1;
    // rom_array[14914] = 32'hFFFFFFF1;
    // rom_array[14915] = 32'hFFFFFFF1;
    // rom_array[14916] = 32'hFFFFFFF1;
    // rom_array[14917] = 32'hFFFFFFF1;
    // rom_array[14918] = 32'hFFFFFFF1;
    // rom_array[14919] = 32'hFFFFFFF1;
    // rom_array[14920] = 32'hFFFFFFF1;
    // rom_array[14921] = 32'hFFFFFFF1;
    // rom_array[14922] = 32'hFFFFFFF1;
    // rom_array[14923] = 32'hFFFFFFF1;
    // rom_array[14924] = 32'hFFFFFFF1;
    // rom_array[14925] = 32'hFFFFFFF1;
    // rom_array[14926] = 32'hFFFFFFF1;
    // rom_array[14927] = 32'hFFFFFFF1;
    // rom_array[14928] = 32'hFFFFFFF1;
    // rom_array[14929] = 32'hFFFFFFF1;
    // rom_array[14930] = 32'hFFFFFFF1;
    // rom_array[14931] = 32'hFFFFFFF1;
    // rom_array[14932] = 32'hFFFFFFF1;
    // rom_array[14933] = 32'hFFFFFFF1;
    // rom_array[14934] = 32'hFFFFFFF1;
    // rom_array[14935] = 32'hFFFFFFF1;
    // rom_array[14936] = 32'hFFFFFFF1;
    // rom_array[14937] = 32'hFFFFFFF1;
    // rom_array[14938] = 32'hFFFFFFF1;
    // rom_array[14939] = 32'hFFFFFFF1;
    // rom_array[14940] = 32'hFFFFFFF1;
    // rom_array[14941] = 32'hFFFFFFF1;
    // rom_array[14942] = 32'hFFFFFFF1;
    // rom_array[14943] = 32'hFFFFFFF1;
    // rom_array[14944] = 32'hFFFFFFF1;
    // rom_array[14945] = 32'hFFFFFFF1;
    // rom_array[14946] = 32'hFFFFFFF1;
    // rom_array[14947] = 32'hFFFFFFF1;
    // rom_array[14948] = 32'hFFFFFFF1;
    // rom_array[14949] = 32'hFFFFFFF1;
    // rom_array[14950] = 32'hFFFFFFF1;
    // rom_array[14951] = 32'hFFFFFFF1;
    // rom_array[14952] = 32'hFFFFFFF1;
    // rom_array[14953] = 32'hFFFFFFF1;
    // rom_array[14954] = 32'hFFFFFFF1;
    // rom_array[14955] = 32'hFFFFFFF1;
    // rom_array[14956] = 32'hFFFFFFF1;
    // rom_array[14957] = 32'hFFFFFFF1;
    // rom_array[14958] = 32'hFFFFFFF1;
    // rom_array[14959] = 32'hFFFFFFF1;
    // rom_array[14960] = 32'hFFFFFFF1;
    // rom_array[14961] = 32'hFFFFFFF1;
    // rom_array[14962] = 32'hFFFFFFF1;
    // rom_array[14963] = 32'hFFFFFFF1;
    // rom_array[14964] = 32'hFFFFFFF1;
    // rom_array[14965] = 32'hFFFFFFF1;
    // rom_array[14966] = 32'hFFFFFFF1;
    // rom_array[14967] = 32'hFFFFFFF1;
    // rom_array[14968] = 32'hFFFFFFF1;
    // rom_array[14969] = 32'hFFFFFFF0;
    // rom_array[14970] = 32'hFFFFFFF0;
    // rom_array[14971] = 32'hFFFFFFF0;
    // rom_array[14972] = 32'hFFFFFFF0;
    // rom_array[14973] = 32'hFFFFFFF0;
    // rom_array[14974] = 32'hFFFFFFF0;
    // rom_array[14975] = 32'hFFFFFFF1;
    // rom_array[14976] = 32'hFFFFFFF1;
    // rom_array[14977] = 32'hFFFFFFF0;
    // rom_array[14978] = 32'hFFFFFFF0;
    // rom_array[14979] = 32'hFFFFFFF0;
    // rom_array[14980] = 32'hFFFFFFF0;
    // rom_array[14981] = 32'hFFFFFFF0;
    // rom_array[14982] = 32'hFFFFFFF0;
    // rom_array[14983] = 32'hFFFFFFF1;
    // rom_array[14984] = 32'hFFFFFFF1;
    // rom_array[14985] = 32'hFFFFFFF0;
    // rom_array[14986] = 32'hFFFFFFF0;
    // rom_array[14987] = 32'hFFFFFFF0;
    // rom_array[14988] = 32'hFFFFFFF0;
    // rom_array[14989] = 32'hFFFFFFF1;
    // rom_array[14990] = 32'hFFFFFFF1;
    // rom_array[14991] = 32'hFFFFFFF1;
    // rom_array[14992] = 32'hFFFFFFF1;
    // rom_array[14993] = 32'hFFFFFFF0;
    // rom_array[14994] = 32'hFFFFFFF0;
    // rom_array[14995] = 32'hFFFFFFF0;
    // rom_array[14996] = 32'hFFFFFFF0;
    // rom_array[14997] = 32'hFFFFFFF1;
    // rom_array[14998] = 32'hFFFFFFF1;
    // rom_array[14999] = 32'hFFFFFFF1;
    // rom_array[15000] = 32'hFFFFFFF1;
    // rom_array[15001] = 32'hFFFFFFF0;
    // rom_array[15002] = 32'hFFFFFFF0;
    // rom_array[15003] = 32'hFFFFFFF1;
    // rom_array[15004] = 32'hFFFFFFF1;
    // rom_array[15005] = 32'hFFFFFFF0;
    // rom_array[15006] = 32'hFFFFFFF0;
    // rom_array[15007] = 32'hFFFFFFF1;
    // rom_array[15008] = 32'hFFFFFFF1;
    // rom_array[15009] = 32'hFFFFFFF0;
    // rom_array[15010] = 32'hFFFFFFF0;
    // rom_array[15011] = 32'hFFFFFFF1;
    // rom_array[15012] = 32'hFFFFFFF1;
    // rom_array[15013] = 32'hFFFFFFF0;
    // rom_array[15014] = 32'hFFFFFFF0;
    // rom_array[15015] = 32'hFFFFFFF1;
    // rom_array[15016] = 32'hFFFFFFF1;
    // rom_array[15017] = 32'hFFFFFFF0;
    // rom_array[15018] = 32'hFFFFFFF0;
    // rom_array[15019] = 32'hFFFFFFF0;
    // rom_array[15020] = 32'hFFFFFFF0;
    // rom_array[15021] = 32'hFFFFFFF1;
    // rom_array[15022] = 32'hFFFFFFF1;
    // rom_array[15023] = 32'hFFFFFFF1;
    // rom_array[15024] = 32'hFFFFFFF1;
    // rom_array[15025] = 32'hFFFFFFF0;
    // rom_array[15026] = 32'hFFFFFFF0;
    // rom_array[15027] = 32'hFFFFFFF0;
    // rom_array[15028] = 32'hFFFFFFF0;
    // rom_array[15029] = 32'hFFFFFFF1;
    // rom_array[15030] = 32'hFFFFFFF1;
    // rom_array[15031] = 32'hFFFFFFF1;
    // rom_array[15032] = 32'hFFFFFFF1;
    // rom_array[15033] = 32'hFFFFFFF0;
    // rom_array[15034] = 32'hFFFFFFF0;
    // rom_array[15035] = 32'hFFFFFFF0;
    // rom_array[15036] = 32'hFFFFFFF0;
    // rom_array[15037] = 32'hFFFFFFF1;
    // rom_array[15038] = 32'hFFFFFFF1;
    // rom_array[15039] = 32'hFFFFFFF1;
    // rom_array[15040] = 32'hFFFFFFF1;
    // rom_array[15041] = 32'hFFFFFFF0;
    // rom_array[15042] = 32'hFFFFFFF0;
    // rom_array[15043] = 32'hFFFFFFF0;
    // rom_array[15044] = 32'hFFFFFFF0;
    // rom_array[15045] = 32'hFFFFFFF1;
    // rom_array[15046] = 32'hFFFFFFF1;
    // rom_array[15047] = 32'hFFFFFFF1;
    // rom_array[15048] = 32'hFFFFFFF1;
    // rom_array[15049] = 32'hFFFFFFF0;
    // rom_array[15050] = 32'hFFFFFFF0;
    // rom_array[15051] = 32'hFFFFFFF1;
    // rom_array[15052] = 32'hFFFFFFF1;
    // rom_array[15053] = 32'hFFFFFFF0;
    // rom_array[15054] = 32'hFFFFFFF0;
    // rom_array[15055] = 32'hFFFFFFF1;
    // rom_array[15056] = 32'hFFFFFFF1;
    // rom_array[15057] = 32'hFFFFFFF0;
    // rom_array[15058] = 32'hFFFFFFF0;
    // rom_array[15059] = 32'hFFFFFFF1;
    // rom_array[15060] = 32'hFFFFFFF1;
    // rom_array[15061] = 32'hFFFFFFF0;
    // rom_array[15062] = 32'hFFFFFFF0;
    // rom_array[15063] = 32'hFFFFFFF1;
    // rom_array[15064] = 32'hFFFFFFF1;
    // rom_array[15065] = 32'hFFFFFFF0;
    // rom_array[15066] = 32'hFFFFFFF0;
    // rom_array[15067] = 32'hFFFFFFF1;
    // rom_array[15068] = 32'hFFFFFFF1;
    // rom_array[15069] = 32'hFFFFFFF0;
    // rom_array[15070] = 32'hFFFFFFF0;
    // rom_array[15071] = 32'hFFFFFFF1;
    // rom_array[15072] = 32'hFFFFFFF1;
    // rom_array[15073] = 32'hFFFFFFF0;
    // rom_array[15074] = 32'hFFFFFFF0;
    // rom_array[15075] = 32'hFFFFFFF1;
    // rom_array[15076] = 32'hFFFFFFF1;
    // rom_array[15077] = 32'hFFFFFFF0;
    // rom_array[15078] = 32'hFFFFFFF0;
    // rom_array[15079] = 32'hFFFFFFF1;
    // rom_array[15080] = 32'hFFFFFFF1;
    // rom_array[15081] = 32'hFFFFFFF0;
    // rom_array[15082] = 32'hFFFFFFF0;
    // rom_array[15083] = 32'hFFFFFFF1;
    // rom_array[15084] = 32'hFFFFFFF1;
    // rom_array[15085] = 32'hFFFFFFF0;
    // rom_array[15086] = 32'hFFFFFFF0;
    // rom_array[15087] = 32'hFFFFFFF0;
    // rom_array[15088] = 32'hFFFFFFF0;
    // rom_array[15089] = 32'hFFFFFFF0;
    // rom_array[15090] = 32'hFFFFFFF0;
    // rom_array[15091] = 32'hFFFFFFF1;
    // rom_array[15092] = 32'hFFFFFFF1;
    // rom_array[15093] = 32'hFFFFFFF0;
    // rom_array[15094] = 32'hFFFFFFF0;
    // rom_array[15095] = 32'hFFFFFFF0;
    // rom_array[15096] = 32'hFFFFFFF0;
    // rom_array[15097] = 32'hFFFFFFF1;
    // rom_array[15098] = 32'hFFFFFFF1;
    // rom_array[15099] = 32'hFFFFFFF1;
    // rom_array[15100] = 32'hFFFFFFF1;
    // rom_array[15101] = 32'hFFFFFFF0;
    // rom_array[15102] = 32'hFFFFFFF0;
    // rom_array[15103] = 32'hFFFFFFF0;
    // rom_array[15104] = 32'hFFFFFFF0;
    // rom_array[15105] = 32'hFFFFFFF1;
    // rom_array[15106] = 32'hFFFFFFF1;
    // rom_array[15107] = 32'hFFFFFFF1;
    // rom_array[15108] = 32'hFFFFFFF1;
    // rom_array[15109] = 32'hFFFFFFF0;
    // rom_array[15110] = 32'hFFFFFFF0;
    // rom_array[15111] = 32'hFFFFFFF0;
    // rom_array[15112] = 32'hFFFFFFF0;
    // rom_array[15113] = 32'hFFFFFFF1;
    // rom_array[15114] = 32'hFFFFFFF1;
    // rom_array[15115] = 32'hFFFFFFF1;
    // rom_array[15116] = 32'hFFFFFFF1;
    // rom_array[15117] = 32'hFFFFFFF0;
    // rom_array[15118] = 32'hFFFFFFF0;
    // rom_array[15119] = 32'hFFFFFFF0;
    // rom_array[15120] = 32'hFFFFFFF0;
    // rom_array[15121] = 32'hFFFFFFF1;
    // rom_array[15122] = 32'hFFFFFFF1;
    // rom_array[15123] = 32'hFFFFFFF1;
    // rom_array[15124] = 32'hFFFFFFF1;
    // rom_array[15125] = 32'hFFFFFFF0;
    // rom_array[15126] = 32'hFFFFFFF0;
    // rom_array[15127] = 32'hFFFFFFF0;
    // rom_array[15128] = 32'hFFFFFFF0;
    // rom_array[15129] = 32'hFFFFFFF1;
    // rom_array[15130] = 32'hFFFFFFF1;
    // rom_array[15131] = 32'hFFFFFFF1;
    // rom_array[15132] = 32'hFFFFFFF1;
    // rom_array[15133] = 32'hFFFFFFF0;
    // rom_array[15134] = 32'hFFFFFFF0;
    // rom_array[15135] = 32'hFFFFFFF0;
    // rom_array[15136] = 32'hFFFFFFF0;
    // rom_array[15137] = 32'hFFFFFFF1;
    // rom_array[15138] = 32'hFFFFFFF1;
    // rom_array[15139] = 32'hFFFFFFF1;
    // rom_array[15140] = 32'hFFFFFFF1;
    // rom_array[15141] = 32'hFFFFFFF0;
    // rom_array[15142] = 32'hFFFFFFF0;
    // rom_array[15143] = 32'hFFFFFFF0;
    // rom_array[15144] = 32'hFFFFFFF0;
    // rom_array[15145] = 32'hFFFFFFF0;
    // rom_array[15146] = 32'hFFFFFFF0;
    // rom_array[15147] = 32'hFFFFFFF0;
    // rom_array[15148] = 32'hFFFFFFF0;
    // rom_array[15149] = 32'hFFFFFFF1;
    // rom_array[15150] = 32'hFFFFFFF1;
    // rom_array[15151] = 32'hFFFFFFF1;
    // rom_array[15152] = 32'hFFFFFFF1;
    // rom_array[15153] = 32'hFFFFFFF0;
    // rom_array[15154] = 32'hFFFFFFF0;
    // rom_array[15155] = 32'hFFFFFFF0;
    // rom_array[15156] = 32'hFFFFFFF0;
    // rom_array[15157] = 32'hFFFFFFF1;
    // rom_array[15158] = 32'hFFFFFFF1;
    // rom_array[15159] = 32'hFFFFFFF1;
    // rom_array[15160] = 32'hFFFFFFF1;
    // rom_array[15161] = 32'hFFFFFFF0;
    // rom_array[15162] = 32'hFFFFFFF0;
    // rom_array[15163] = 32'hFFFFFFF0;
    // rom_array[15164] = 32'hFFFFFFF0;
    // rom_array[15165] = 32'hFFFFFFF1;
    // rom_array[15166] = 32'hFFFFFFF1;
    // rom_array[15167] = 32'hFFFFFFF1;
    // rom_array[15168] = 32'hFFFFFFF1;
    // rom_array[15169] = 32'hFFFFFFF0;
    // rom_array[15170] = 32'hFFFFFFF0;
    // rom_array[15171] = 32'hFFFFFFF0;
    // rom_array[15172] = 32'hFFFFFFF0;
    // rom_array[15173] = 32'hFFFFFFF1;
    // rom_array[15174] = 32'hFFFFFFF1;
    // rom_array[15175] = 32'hFFFFFFF1;
    // rom_array[15176] = 32'hFFFFFFF1;
    // rom_array[15177] = 32'hFFFFFFF0;
    // rom_array[15178] = 32'hFFFFFFF0;
    // rom_array[15179] = 32'hFFFFFFF0;
    // rom_array[15180] = 32'hFFFFFFF0;
    // rom_array[15181] = 32'hFFFFFFF1;
    // rom_array[15182] = 32'hFFFFFFF1;
    // rom_array[15183] = 32'hFFFFFFF1;
    // rom_array[15184] = 32'hFFFFFFF1;
    // rom_array[15185] = 32'hFFFFFFF0;
    // rom_array[15186] = 32'hFFFFFFF0;
    // rom_array[15187] = 32'hFFFFFFF0;
    // rom_array[15188] = 32'hFFFFFFF0;
    // rom_array[15189] = 32'hFFFFFFF1;
    // rom_array[15190] = 32'hFFFFFFF1;
    // rom_array[15191] = 32'hFFFFFFF1;
    // rom_array[15192] = 32'hFFFFFFF1;
    // rom_array[15193] = 32'hFFFFFFF1;
    // rom_array[15194] = 32'hFFFFFFF1;
    // rom_array[15195] = 32'hFFFFFFF1;
    // rom_array[15196] = 32'hFFFFFFF1;
    // rom_array[15197] = 32'hFFFFFFF1;
    // rom_array[15198] = 32'hFFFFFFF1;
    // rom_array[15199] = 32'hFFFFFFF1;
    // rom_array[15200] = 32'hFFFFFFF1;
    // rom_array[15201] = 32'hFFFFFFF1;
    // rom_array[15202] = 32'hFFFFFFF1;
    // rom_array[15203] = 32'hFFFFFFF1;
    // rom_array[15204] = 32'hFFFFFFF1;
    // rom_array[15205] = 32'hFFFFFFF1;
    // rom_array[15206] = 32'hFFFFFFF1;
    // rom_array[15207] = 32'hFFFFFFF1;
    // rom_array[15208] = 32'hFFFFFFF1;
    // rom_array[15209] = 32'hFFFFFFF1;
    // rom_array[15210] = 32'hFFFFFFF1;
    // rom_array[15211] = 32'hFFFFFFF1;
    // rom_array[15212] = 32'hFFFFFFF1;
    // rom_array[15213] = 32'hFFFFFFF1;
    // rom_array[15214] = 32'hFFFFFFF1;
    // rom_array[15215] = 32'hFFFFFFF1;
    // rom_array[15216] = 32'hFFFFFFF1;
    // rom_array[15217] = 32'hFFFFFFF1;
    // rom_array[15218] = 32'hFFFFFFF1;
    // rom_array[15219] = 32'hFFFFFFF1;
    // rom_array[15220] = 32'hFFFFFFF1;
    // rom_array[15221] = 32'hFFFFFFF1;
    // rom_array[15222] = 32'hFFFFFFF1;
    // rom_array[15223] = 32'hFFFFFFF1;
    // rom_array[15224] = 32'hFFFFFFF1;
    // rom_array[15225] = 32'hFFFFFFF1;
    // rom_array[15226] = 32'hFFFFFFF1;
    // rom_array[15227] = 32'hFFFFFFF1;
    // rom_array[15228] = 32'hFFFFFFF1;
    // rom_array[15229] = 32'hFFFFFFF1;
    // rom_array[15230] = 32'hFFFFFFF1;
    // rom_array[15231] = 32'hFFFFFFF1;
    // rom_array[15232] = 32'hFFFFFFF1;
    // rom_array[15233] = 32'hFFFFFFF1;
    // rom_array[15234] = 32'hFFFFFFF1;
    // rom_array[15235] = 32'hFFFFFFF1;
    // rom_array[15236] = 32'hFFFFFFF1;
    // rom_array[15237] = 32'hFFFFFFF1;
    // rom_array[15238] = 32'hFFFFFFF1;
    // rom_array[15239] = 32'hFFFFFFF1;
    // rom_array[15240] = 32'hFFFFFFF1;
    // rom_array[15241] = 32'hFFFFFFF1;
    // rom_array[15242] = 32'hFFFFFFF1;
    // rom_array[15243] = 32'hFFFFFFF1;
    // rom_array[15244] = 32'hFFFFFFF1;
    // rom_array[15245] = 32'hFFFFFFF1;
    // rom_array[15246] = 32'hFFFFFFF1;
    // rom_array[15247] = 32'hFFFFFFF1;
    // rom_array[15248] = 32'hFFFFFFF1;
    // rom_array[15249] = 32'hFFFFFFF1;
    // rom_array[15250] = 32'hFFFFFFF1;
    // rom_array[15251] = 32'hFFFFFFF1;
    // rom_array[15252] = 32'hFFFFFFF1;
    // rom_array[15253] = 32'hFFFFFFF1;
    // rom_array[15254] = 32'hFFFFFFF1;
    // rom_array[15255] = 32'hFFFFFFF1;
    // rom_array[15256] = 32'hFFFFFFF1;
    // rom_array[15257] = 32'hFFFFFFF0;
    // rom_array[15258] = 32'hFFFFFFF0;
    // rom_array[15259] = 32'hFFFFFFF0;
    // rom_array[15260] = 32'hFFFFFFF0;
    // rom_array[15261] = 32'hFFFFFFF1;
    // rom_array[15262] = 32'hFFFFFFF1;
    // rom_array[15263] = 32'hFFFFFFF1;
    // rom_array[15264] = 32'hFFFFFFF1;
    // rom_array[15265] = 32'hFFFFFFF0;
    // rom_array[15266] = 32'hFFFFFFF0;
    // rom_array[15267] = 32'hFFFFFFF0;
    // rom_array[15268] = 32'hFFFFFFF0;
    // rom_array[15269] = 32'hFFFFFFF1;
    // rom_array[15270] = 32'hFFFFFFF1;
    // rom_array[15271] = 32'hFFFFFFF1;
    // rom_array[15272] = 32'hFFFFFFF1;
    // rom_array[15273] = 32'hFFFFFFF0;
    // rom_array[15274] = 32'hFFFFFFF0;
    // rom_array[15275] = 32'hFFFFFFF0;
    // rom_array[15276] = 32'hFFFFFFF0;
    // rom_array[15277] = 32'hFFFFFFF1;
    // rom_array[15278] = 32'hFFFFFFF1;
    // rom_array[15279] = 32'hFFFFFFF1;
    // rom_array[15280] = 32'hFFFFFFF1;
    // rom_array[15281] = 32'hFFFFFFF0;
    // rom_array[15282] = 32'hFFFFFFF0;
    // rom_array[15283] = 32'hFFFFFFF0;
    // rom_array[15284] = 32'hFFFFFFF0;
    // rom_array[15285] = 32'hFFFFFFF1;
    // rom_array[15286] = 32'hFFFFFFF1;
    // rom_array[15287] = 32'hFFFFFFF1;
    // rom_array[15288] = 32'hFFFFFFF1;
    // rom_array[15289] = 32'hFFFFFFF0;
    // rom_array[15290] = 32'hFFFFFFF0;
    // rom_array[15291] = 32'hFFFFFFF0;
    // rom_array[15292] = 32'hFFFFFFF0;
    // rom_array[15293] = 32'hFFFFFFF1;
    // rom_array[15294] = 32'hFFFFFFF1;
    // rom_array[15295] = 32'hFFFFFFF1;
    // rom_array[15296] = 32'hFFFFFFF1;
    // rom_array[15297] = 32'hFFFFFFF0;
    // rom_array[15298] = 32'hFFFFFFF0;
    // rom_array[15299] = 32'hFFFFFFF0;
    // rom_array[15300] = 32'hFFFFFFF0;
    // rom_array[15301] = 32'hFFFFFFF1;
    // rom_array[15302] = 32'hFFFFFFF1;
    // rom_array[15303] = 32'hFFFFFFF1;
    // rom_array[15304] = 32'hFFFFFFF1;
    // rom_array[15305] = 32'hFFFFFFF0;
    // rom_array[15306] = 32'hFFFFFFF0;
    // rom_array[15307] = 32'hFFFFFFF0;
    // rom_array[15308] = 32'hFFFFFFF0;
    // rom_array[15309] = 32'hFFFFFFF1;
    // rom_array[15310] = 32'hFFFFFFF1;
    // rom_array[15311] = 32'hFFFFFFF1;
    // rom_array[15312] = 32'hFFFFFFF1;
    // rom_array[15313] = 32'hFFFFFFF0;
    // rom_array[15314] = 32'hFFFFFFF0;
    // rom_array[15315] = 32'hFFFFFFF0;
    // rom_array[15316] = 32'hFFFFFFF0;
    // rom_array[15317] = 32'hFFFFFFF1;
    // rom_array[15318] = 32'hFFFFFFF1;
    // rom_array[15319] = 32'hFFFFFFF1;
    // rom_array[15320] = 32'hFFFFFFF1;
    // rom_array[15321] = 32'hFFFFFFF1;
    // rom_array[15322] = 32'hFFFFFFF1;
    // rom_array[15323] = 32'hFFFFFFF1;
    // rom_array[15324] = 32'hFFFFFFF1;
    // rom_array[15325] = 32'hFFFFFFF1;
    // rom_array[15326] = 32'hFFFFFFF1;
    // rom_array[15327] = 32'hFFFFFFF1;
    // rom_array[15328] = 32'hFFFFFFF1;
    // rom_array[15329] = 32'hFFFFFFF1;
    // rom_array[15330] = 32'hFFFFFFF1;
    // rom_array[15331] = 32'hFFFFFFF1;
    // rom_array[15332] = 32'hFFFFFFF1;
    // rom_array[15333] = 32'hFFFFFFF1;
    // rom_array[15334] = 32'hFFFFFFF1;
    // rom_array[15335] = 32'hFFFFFFF1;
    // rom_array[15336] = 32'hFFFFFFF1;
    // rom_array[15337] = 32'hFFFFFFF1;
    // rom_array[15338] = 32'hFFFFFFF1;
    // rom_array[15339] = 32'hFFFFFFF1;
    // rom_array[15340] = 32'hFFFFFFF1;
    // rom_array[15341] = 32'hFFFFFFF1;
    // rom_array[15342] = 32'hFFFFFFF1;
    // rom_array[15343] = 32'hFFFFFFF1;
    // rom_array[15344] = 32'hFFFFFFF1;
    // rom_array[15345] = 32'hFFFFFFF1;
    // rom_array[15346] = 32'hFFFFFFF1;
    // rom_array[15347] = 32'hFFFFFFF1;
    // rom_array[15348] = 32'hFFFFFFF1;
    // rom_array[15349] = 32'hFFFFFFF1;
    // rom_array[15350] = 32'hFFFFFFF1;
    // rom_array[15351] = 32'hFFFFFFF1;
    // rom_array[15352] = 32'hFFFFFFF1;
    // rom_array[15353] = 32'hFFFFFFF1;
    // rom_array[15354] = 32'hFFFFFFF1;
    // rom_array[15355] = 32'hFFFFFFF1;
    // rom_array[15356] = 32'hFFFFFFF1;
    // rom_array[15357] = 32'hFFFFFFF1;
    // rom_array[15358] = 32'hFFFFFFF1;
    // rom_array[15359] = 32'hFFFFFFF1;
    // rom_array[15360] = 32'hFFFFFFF1;
    // rom_array[15361] = 32'hFFFFFFF1;
    // rom_array[15362] = 32'hFFFFFFF1;
    // rom_array[15363] = 32'hFFFFFFF1;
    // rom_array[15364] = 32'hFFFFFFF1;
    // rom_array[15365] = 32'hFFFFFFF1;
    // rom_array[15366] = 32'hFFFFFFF1;
    // rom_array[15367] = 32'hFFFFFFF1;
    // rom_array[15368] = 32'hFFFFFFF1;
    // rom_array[15369] = 32'hFFFFFFF1;
    // rom_array[15370] = 32'hFFFFFFF1;
    // rom_array[15371] = 32'hFFFFFFF1;
    // rom_array[15372] = 32'hFFFFFFF1;
    // rom_array[15373] = 32'hFFFFFFF1;
    // rom_array[15374] = 32'hFFFFFFF1;
    // rom_array[15375] = 32'hFFFFFFF1;
    // rom_array[15376] = 32'hFFFFFFF1;
    // rom_array[15377] = 32'hFFFFFFF1;
    // rom_array[15378] = 32'hFFFFFFF1;
    // rom_array[15379] = 32'hFFFFFFF1;
    // rom_array[15380] = 32'hFFFFFFF1;
    // rom_array[15381] = 32'hFFFFFFF1;
    // rom_array[15382] = 32'hFFFFFFF1;
    // rom_array[15383] = 32'hFFFFFFF1;
    // rom_array[15384] = 32'hFFFFFFF1;
    // rom_array[15385] = 32'hFFFFFFF1;
    // rom_array[15386] = 32'hFFFFFFF1;
    // rom_array[15387] = 32'hFFFFFFF1;
    // rom_array[15388] = 32'hFFFFFFF1;
    // rom_array[15389] = 32'hFFFFFFF0;
    // rom_array[15390] = 32'hFFFFFFF0;
    // rom_array[15391] = 32'hFFFFFFF0;
    // rom_array[15392] = 32'hFFFFFFF0;
    // rom_array[15393] = 32'hFFFFFFF1;
    // rom_array[15394] = 32'hFFFFFFF1;
    // rom_array[15395] = 32'hFFFFFFF1;
    // rom_array[15396] = 32'hFFFFFFF1;
    // rom_array[15397] = 32'hFFFFFFF0;
    // rom_array[15398] = 32'hFFFFFFF0;
    // rom_array[15399] = 32'hFFFFFFF0;
    // rom_array[15400] = 32'hFFFFFFF0;
    // rom_array[15401] = 32'hFFFFFFF1;
    // rom_array[15402] = 32'hFFFFFFF1;
    // rom_array[15403] = 32'hFFFFFFF1;
    // rom_array[15404] = 32'hFFFFFFF1;
    // rom_array[15405] = 32'hFFFFFFF0;
    // rom_array[15406] = 32'hFFFFFFF0;
    // rom_array[15407] = 32'hFFFFFFF0;
    // rom_array[15408] = 32'hFFFFFFF0;
    // rom_array[15409] = 32'hFFFFFFF1;
    // rom_array[15410] = 32'hFFFFFFF1;
    // rom_array[15411] = 32'hFFFFFFF1;
    // rom_array[15412] = 32'hFFFFFFF1;
    // rom_array[15413] = 32'hFFFFFFF0;
    // rom_array[15414] = 32'hFFFFFFF0;
    // rom_array[15415] = 32'hFFFFFFF0;
    // rom_array[15416] = 32'hFFFFFFF0;
    // rom_array[15417] = 32'hFFFFFFF1;
    // rom_array[15418] = 32'hFFFFFFF1;
    // rom_array[15419] = 32'hFFFFFFF1;
    // rom_array[15420] = 32'hFFFFFFF1;
    // rom_array[15421] = 32'hFFFFFFF0;
    // rom_array[15422] = 32'hFFFFFFF0;
    // rom_array[15423] = 32'hFFFFFFF0;
    // rom_array[15424] = 32'hFFFFFFF0;
    // rom_array[15425] = 32'hFFFFFFF1;
    // rom_array[15426] = 32'hFFFFFFF1;
    // rom_array[15427] = 32'hFFFFFFF1;
    // rom_array[15428] = 32'hFFFFFFF1;
    // rom_array[15429] = 32'hFFFFFFF0;
    // rom_array[15430] = 32'hFFFFFFF0;
    // rom_array[15431] = 32'hFFFFFFF0;
    // rom_array[15432] = 32'hFFFFFFF0;
    // rom_array[15433] = 32'hFFFFFFF1;
    // rom_array[15434] = 32'hFFFFFFF1;
    // rom_array[15435] = 32'hFFFFFFF1;
    // rom_array[15436] = 32'hFFFFFFF1;
    // rom_array[15437] = 32'hFFFFFFF0;
    // rom_array[15438] = 32'hFFFFFFF0;
    // rom_array[15439] = 32'hFFFFFFF0;
    // rom_array[15440] = 32'hFFFFFFF0;
    // rom_array[15441] = 32'hFFFFFFF1;
    // rom_array[15442] = 32'hFFFFFFF1;
    // rom_array[15443] = 32'hFFFFFFF1;
    // rom_array[15444] = 32'hFFFFFFF1;
    // rom_array[15445] = 32'hFFFFFFF0;
    // rom_array[15446] = 32'hFFFFFFF0;
    // rom_array[15447] = 32'hFFFFFFF0;
    // rom_array[15448] = 32'hFFFFFFF0;
    // rom_array[15449] = 32'hFFFFFFF1;
    // rom_array[15450] = 32'hFFFFFFF1;
    // rom_array[15451] = 32'hFFFFFFF1;
    // rom_array[15452] = 32'hFFFFFFF1;
    // rom_array[15453] = 32'hFFFFFFF0;
    // rom_array[15454] = 32'hFFFFFFF0;
    // rom_array[15455] = 32'hFFFFFFF0;
    // rom_array[15456] = 32'hFFFFFFF0;
    // rom_array[15457] = 32'hFFFFFFF1;
    // rom_array[15458] = 32'hFFFFFFF1;
    // rom_array[15459] = 32'hFFFFFFF1;
    // rom_array[15460] = 32'hFFFFFFF1;
    // rom_array[15461] = 32'hFFFFFFF0;
    // rom_array[15462] = 32'hFFFFFFF0;
    // rom_array[15463] = 32'hFFFFFFF0;
    // rom_array[15464] = 32'hFFFFFFF0;
    // rom_array[15465] = 32'hFFFFFFF1;
    // rom_array[15466] = 32'hFFFFFFF1;
    // rom_array[15467] = 32'hFFFFFFF1;
    // rom_array[15468] = 32'hFFFFFFF1;
    // rom_array[15469] = 32'hFFFFFFF0;
    // rom_array[15470] = 32'hFFFFFFF0;
    // rom_array[15471] = 32'hFFFFFFF0;
    // rom_array[15472] = 32'hFFFFFFF0;
    // rom_array[15473] = 32'hFFFFFFF1;
    // rom_array[15474] = 32'hFFFFFFF1;
    // rom_array[15475] = 32'hFFFFFFF1;
    // rom_array[15476] = 32'hFFFFFFF1;
    // rom_array[15477] = 32'hFFFFFFF0;
    // rom_array[15478] = 32'hFFFFFFF0;
    // rom_array[15479] = 32'hFFFFFFF0;
    // rom_array[15480] = 32'hFFFFFFF0;
    // rom_array[15481] = 32'hFFFFFFF1;
    // rom_array[15482] = 32'hFFFFFFF1;
    // rom_array[15483] = 32'hFFFFFFF1;
    // rom_array[15484] = 32'hFFFFFFF1;
    // rom_array[15485] = 32'hFFFFFFF0;
    // rom_array[15486] = 32'hFFFFFFF0;
    // rom_array[15487] = 32'hFFFFFFF0;
    // rom_array[15488] = 32'hFFFFFFF0;
    // rom_array[15489] = 32'hFFFFFFF1;
    // rom_array[15490] = 32'hFFFFFFF1;
    // rom_array[15491] = 32'hFFFFFFF1;
    // rom_array[15492] = 32'hFFFFFFF1;
    // rom_array[15493] = 32'hFFFFFFF0;
    // rom_array[15494] = 32'hFFFFFFF0;
    // rom_array[15495] = 32'hFFFFFFF0;
    // rom_array[15496] = 32'hFFFFFFF0;
    // rom_array[15497] = 32'hFFFFFFF1;
    // rom_array[15498] = 32'hFFFFFFF1;
    // rom_array[15499] = 32'hFFFFFFF1;
    // rom_array[15500] = 32'hFFFFFFF1;
    // rom_array[15501] = 32'hFFFFFFF0;
    // rom_array[15502] = 32'hFFFFFFF0;
    // rom_array[15503] = 32'hFFFFFFF0;
    // rom_array[15504] = 32'hFFFFFFF0;
    // rom_array[15505] = 32'hFFFFFFF1;
    // rom_array[15506] = 32'hFFFFFFF1;
    // rom_array[15507] = 32'hFFFFFFF1;
    // rom_array[15508] = 32'hFFFFFFF1;
    // rom_array[15509] = 32'hFFFFFFF0;
    // rom_array[15510] = 32'hFFFFFFF0;
    // rom_array[15511] = 32'hFFFFFFF0;
    // rom_array[15512] = 32'hFFFFFFF0;
    // rom_array[15513] = 32'hFFFFFFF0;
    // rom_array[15514] = 32'hFFFFFFF0;
    // rom_array[15515] = 32'hFFFFFFF0;
    // rom_array[15516] = 32'hFFFFFFF0;
    // rom_array[15517] = 32'hFFFFFFF0;
    // rom_array[15518] = 32'hFFFFFFF0;
    // rom_array[15519] = 32'hFFFFFFF1;
    // rom_array[15520] = 32'hFFFFFFF1;
    // rom_array[15521] = 32'hFFFFFFF0;
    // rom_array[15522] = 32'hFFFFFFF0;
    // rom_array[15523] = 32'hFFFFFFF0;
    // rom_array[15524] = 32'hFFFFFFF0;
    // rom_array[15525] = 32'hFFFFFFF0;
    // rom_array[15526] = 32'hFFFFFFF0;
    // rom_array[15527] = 32'hFFFFFFF1;
    // rom_array[15528] = 32'hFFFFFFF1;
    // rom_array[15529] = 32'hFFFFFFF0;
    // rom_array[15530] = 32'hFFFFFFF0;
    // rom_array[15531] = 32'hFFFFFFF0;
    // rom_array[15532] = 32'hFFFFFFF0;
    // rom_array[15533] = 32'hFFFFFFF1;
    // rom_array[15534] = 32'hFFFFFFF1;
    // rom_array[15535] = 32'hFFFFFFF1;
    // rom_array[15536] = 32'hFFFFFFF1;
    // rom_array[15537] = 32'hFFFFFFF0;
    // rom_array[15538] = 32'hFFFFFFF0;
    // rom_array[15539] = 32'hFFFFFFF0;
    // rom_array[15540] = 32'hFFFFFFF0;
    // rom_array[15541] = 32'hFFFFFFF1;
    // rom_array[15542] = 32'hFFFFFFF1;
    // rom_array[15543] = 32'hFFFFFFF1;
    // rom_array[15544] = 32'hFFFFFFF1;
    // rom_array[15545] = 32'hFFFFFFF0;
    // rom_array[15546] = 32'hFFFFFFF0;
    // rom_array[15547] = 32'hFFFFFFF1;
    // rom_array[15548] = 32'hFFFFFFF1;
    // rom_array[15549] = 32'hFFFFFFF0;
    // rom_array[15550] = 32'hFFFFFFF0;
    // rom_array[15551] = 32'hFFFFFFF1;
    // rom_array[15552] = 32'hFFFFFFF1;
    // rom_array[15553] = 32'hFFFFFFF0;
    // rom_array[15554] = 32'hFFFFFFF0;
    // rom_array[15555] = 32'hFFFFFFF1;
    // rom_array[15556] = 32'hFFFFFFF1;
    // rom_array[15557] = 32'hFFFFFFF0;
    // rom_array[15558] = 32'hFFFFFFF0;
    // rom_array[15559] = 32'hFFFFFFF1;
    // rom_array[15560] = 32'hFFFFFFF1;
    // rom_array[15561] = 32'hFFFFFFF0;
    // rom_array[15562] = 32'hFFFFFFF0;
    // rom_array[15563] = 32'hFFFFFFF0;
    // rom_array[15564] = 32'hFFFFFFF0;
    // rom_array[15565] = 32'hFFFFFFF1;
    // rom_array[15566] = 32'hFFFFFFF1;
    // rom_array[15567] = 32'hFFFFFFF1;
    // rom_array[15568] = 32'hFFFFFFF1;
    // rom_array[15569] = 32'hFFFFFFF0;
    // rom_array[15570] = 32'hFFFFFFF0;
    // rom_array[15571] = 32'hFFFFFFF0;
    // rom_array[15572] = 32'hFFFFFFF0;
    // rom_array[15573] = 32'hFFFFFFF1;
    // rom_array[15574] = 32'hFFFFFFF1;
    // rom_array[15575] = 32'hFFFFFFF1;
    // rom_array[15576] = 32'hFFFFFFF1;
    // rom_array[15577] = 32'hFFFFFFF0;
    // rom_array[15578] = 32'hFFFFFFF0;
    // rom_array[15579] = 32'hFFFFFFF0;
    // rom_array[15580] = 32'hFFFFFFF0;
    // rom_array[15581] = 32'hFFFFFFF1;
    // rom_array[15582] = 32'hFFFFFFF1;
    // rom_array[15583] = 32'hFFFFFFF1;
    // rom_array[15584] = 32'hFFFFFFF1;
    // rom_array[15585] = 32'hFFFFFFF0;
    // rom_array[15586] = 32'hFFFFFFF0;
    // rom_array[15587] = 32'hFFFFFFF0;
    // rom_array[15588] = 32'hFFFFFFF0;
    // rom_array[15589] = 32'hFFFFFFF1;
    // rom_array[15590] = 32'hFFFFFFF1;
    // rom_array[15591] = 32'hFFFFFFF1;
    // rom_array[15592] = 32'hFFFFFFF1;
    // rom_array[15593] = 32'hFFFFFFF0;
    // rom_array[15594] = 32'hFFFFFFF0;
    // rom_array[15595] = 32'hFFFFFFF1;
    // rom_array[15596] = 32'hFFFFFFF1;
    // rom_array[15597] = 32'hFFFFFFF0;
    // rom_array[15598] = 32'hFFFFFFF0;
    // rom_array[15599] = 32'hFFFFFFF1;
    // rom_array[15600] = 32'hFFFFFFF1;
    // rom_array[15601] = 32'hFFFFFFF0;
    // rom_array[15602] = 32'hFFFFFFF0;
    // rom_array[15603] = 32'hFFFFFFF1;
    // rom_array[15604] = 32'hFFFFFFF1;
    // rom_array[15605] = 32'hFFFFFFF0;
    // rom_array[15606] = 32'hFFFFFFF0;
    // rom_array[15607] = 32'hFFFFFFF1;
    // rom_array[15608] = 32'hFFFFFFF1;
    // rom_array[15609] = 32'hFFFFFFF0;
    // rom_array[15610] = 32'hFFFFFFF0;
    // rom_array[15611] = 32'hFFFFFFF1;
    // rom_array[15612] = 32'hFFFFFFF1;
    // rom_array[15613] = 32'hFFFFFFF0;
    // rom_array[15614] = 32'hFFFFFFF0;
    // rom_array[15615] = 32'hFFFFFFF1;
    // rom_array[15616] = 32'hFFFFFFF1;
    // rom_array[15617] = 32'hFFFFFFF0;
    // rom_array[15618] = 32'hFFFFFFF0;
    // rom_array[15619] = 32'hFFFFFFF1;
    // rom_array[15620] = 32'hFFFFFFF1;
    // rom_array[15621] = 32'hFFFFFFF0;
    // rom_array[15622] = 32'hFFFFFFF0;
    // rom_array[15623] = 32'hFFFFFFF1;
    // rom_array[15624] = 32'hFFFFFFF1;
    // rom_array[15625] = 32'hFFFFFFF0;
    // rom_array[15626] = 32'hFFFFFFF0;
    // rom_array[15627] = 32'hFFFFFFF1;
    // rom_array[15628] = 32'hFFFFFFF1;
    // rom_array[15629] = 32'hFFFFFFF0;
    // rom_array[15630] = 32'hFFFFFFF0;
    // rom_array[15631] = 32'hFFFFFFF0;
    // rom_array[15632] = 32'hFFFFFFF0;
    // rom_array[15633] = 32'hFFFFFFF0;
    // rom_array[15634] = 32'hFFFFFFF0;
    // rom_array[15635] = 32'hFFFFFFF1;
    // rom_array[15636] = 32'hFFFFFFF1;
    // rom_array[15637] = 32'hFFFFFFF0;
    // rom_array[15638] = 32'hFFFFFFF0;
    // rom_array[15639] = 32'hFFFFFFF0;
    // rom_array[15640] = 32'hFFFFFFF0;
    // rom_array[15641] = 32'hFFFFFFF1;
    // rom_array[15642] = 32'hFFFFFFF1;
    // rom_array[15643] = 32'hFFFFFFF1;
    // rom_array[15644] = 32'hFFFFFFF1;
    // rom_array[15645] = 32'hFFFFFFF0;
    // rom_array[15646] = 32'hFFFFFFF0;
    // rom_array[15647] = 32'hFFFFFFF0;
    // rom_array[15648] = 32'hFFFFFFF0;
    // rom_array[15649] = 32'hFFFFFFF1;
    // rom_array[15650] = 32'hFFFFFFF1;
    // rom_array[15651] = 32'hFFFFFFF1;
    // rom_array[15652] = 32'hFFFFFFF1;
    // rom_array[15653] = 32'hFFFFFFF0;
    // rom_array[15654] = 32'hFFFFFFF0;
    // rom_array[15655] = 32'hFFFFFFF0;
    // rom_array[15656] = 32'hFFFFFFF0;
    // rom_array[15657] = 32'hFFFFFFF1;
    // rom_array[15658] = 32'hFFFFFFF1;
    // rom_array[15659] = 32'hFFFFFFF1;
    // rom_array[15660] = 32'hFFFFFFF1;
    // rom_array[15661] = 32'hFFFFFFF0;
    // rom_array[15662] = 32'hFFFFFFF0;
    // rom_array[15663] = 32'hFFFFFFF0;
    // rom_array[15664] = 32'hFFFFFFF0;
    // rom_array[15665] = 32'hFFFFFFF1;
    // rom_array[15666] = 32'hFFFFFFF1;
    // rom_array[15667] = 32'hFFFFFFF1;
    // rom_array[15668] = 32'hFFFFFFF1;
    // rom_array[15669] = 32'hFFFFFFF0;
    // rom_array[15670] = 32'hFFFFFFF0;
    // rom_array[15671] = 32'hFFFFFFF0;
    // rom_array[15672] = 32'hFFFFFFF0;
    // rom_array[15673] = 32'hFFFFFFF1;
    // rom_array[15674] = 32'hFFFFFFF1;
    // rom_array[15675] = 32'hFFFFFFF1;
    // rom_array[15676] = 32'hFFFFFFF1;
    // rom_array[15677] = 32'hFFFFFFF0;
    // rom_array[15678] = 32'hFFFFFFF0;
    // rom_array[15679] = 32'hFFFFFFF0;
    // rom_array[15680] = 32'hFFFFFFF0;
    // rom_array[15681] = 32'hFFFFFFF1;
    // rom_array[15682] = 32'hFFFFFFF1;
    // rom_array[15683] = 32'hFFFFFFF1;
    // rom_array[15684] = 32'hFFFFFFF1;
    // rom_array[15685] = 32'hFFFFFFF0;
    // rom_array[15686] = 32'hFFFFFFF0;
    // rom_array[15687] = 32'hFFFFFFF0;
    // rom_array[15688] = 32'hFFFFFFF0;
    // rom_array[15689] = 32'hFFFFFFF0;
    // rom_array[15690] = 32'hFFFFFFF0;
    // rom_array[15691] = 32'hFFFFFFF0;
    // rom_array[15692] = 32'hFFFFFFF0;
    // rom_array[15693] = 32'hFFFFFFF1;
    // rom_array[15694] = 32'hFFFFFFF1;
    // rom_array[15695] = 32'hFFFFFFF1;
    // rom_array[15696] = 32'hFFFFFFF1;
    // rom_array[15697] = 32'hFFFFFFF0;
    // rom_array[15698] = 32'hFFFFFFF0;
    // rom_array[15699] = 32'hFFFFFFF0;
    // rom_array[15700] = 32'hFFFFFFF0;
    // rom_array[15701] = 32'hFFFFFFF1;
    // rom_array[15702] = 32'hFFFFFFF1;
    // rom_array[15703] = 32'hFFFFFFF1;
    // rom_array[15704] = 32'hFFFFFFF1;
    // rom_array[15705] = 32'hFFFFFFF0;
    // rom_array[15706] = 32'hFFFFFFF0;
    // rom_array[15707] = 32'hFFFFFFF0;
    // rom_array[15708] = 32'hFFFFFFF0;
    // rom_array[15709] = 32'hFFFFFFF1;
    // rom_array[15710] = 32'hFFFFFFF1;
    // rom_array[15711] = 32'hFFFFFFF1;
    // rom_array[15712] = 32'hFFFFFFF1;
    // rom_array[15713] = 32'hFFFFFFF0;
    // rom_array[15714] = 32'hFFFFFFF0;
    // rom_array[15715] = 32'hFFFFFFF0;
    // rom_array[15716] = 32'hFFFFFFF0;
    // rom_array[15717] = 32'hFFFFFFF1;
    // rom_array[15718] = 32'hFFFFFFF1;
    // rom_array[15719] = 32'hFFFFFFF1;
    // rom_array[15720] = 32'hFFFFFFF1;
    // rom_array[15721] = 32'hFFFFFFF0;
    // rom_array[15722] = 32'hFFFFFFF0;
    // rom_array[15723] = 32'hFFFFFFF0;
    // rom_array[15724] = 32'hFFFFFFF0;
    // rom_array[15725] = 32'hFFFFFFF1;
    // rom_array[15726] = 32'hFFFFFFF1;
    // rom_array[15727] = 32'hFFFFFFF1;
    // rom_array[15728] = 32'hFFFFFFF1;
    // rom_array[15729] = 32'hFFFFFFF0;
    // rom_array[15730] = 32'hFFFFFFF0;
    // rom_array[15731] = 32'hFFFFFFF0;
    // rom_array[15732] = 32'hFFFFFFF0;
    // rom_array[15733] = 32'hFFFFFFF1;
    // rom_array[15734] = 32'hFFFFFFF1;
    // rom_array[15735] = 32'hFFFFFFF1;
    // rom_array[15736] = 32'hFFFFFFF1;
    // rom_array[15737] = 32'hFFFFFFF0;
    // rom_array[15738] = 32'hFFFFFFF0;
    // rom_array[15739] = 32'hFFFFFFF0;
    // rom_array[15740] = 32'hFFFFFFF0;
    // rom_array[15741] = 32'hFFFFFFF1;
    // rom_array[15742] = 32'hFFFFFFF1;
    // rom_array[15743] = 32'hFFFFFFF1;
    // rom_array[15744] = 32'hFFFFFFF1;
    // rom_array[15745] = 32'hFFFFFFF0;
    // rom_array[15746] = 32'hFFFFFFF0;
    // rom_array[15747] = 32'hFFFFFFF0;
    // rom_array[15748] = 32'hFFFFFFF0;
    // rom_array[15749] = 32'hFFFFFFF1;
    // rom_array[15750] = 32'hFFFFFFF1;
    // rom_array[15751] = 32'hFFFFFFF1;
    // rom_array[15752] = 32'hFFFFFFF1;
    // rom_array[15753] = 32'hFFFFFFF0;
    // rom_array[15754] = 32'hFFFFFFF0;
    // rom_array[15755] = 32'hFFFFFFF0;
    // rom_array[15756] = 32'hFFFFFFF0;
    // rom_array[15757] = 32'hFFFFFFF1;
    // rom_array[15758] = 32'hFFFFFFF1;
    // rom_array[15759] = 32'hFFFFFFF1;
    // rom_array[15760] = 32'hFFFFFFF1;
    // rom_array[15761] = 32'hFFFFFFF0;
    // rom_array[15762] = 32'hFFFFFFF0;
    // rom_array[15763] = 32'hFFFFFFF0;
    // rom_array[15764] = 32'hFFFFFFF0;
    // rom_array[15765] = 32'hFFFFFFF1;
    // rom_array[15766] = 32'hFFFFFFF1;
    // rom_array[15767] = 32'hFFFFFFF1;
    // rom_array[15768] = 32'hFFFFFFF1;
    // rom_array[15769] = 32'hFFFFFFF0;
    // rom_array[15770] = 32'hFFFFFFF0;
    // rom_array[15771] = 32'hFFFFFFF0;
    // rom_array[15772] = 32'hFFFFFFF0;
    // rom_array[15773] = 32'hFFFFFFF1;
    // rom_array[15774] = 32'hFFFFFFF1;
    // rom_array[15775] = 32'hFFFFFFF1;
    // rom_array[15776] = 32'hFFFFFFF1;
    // rom_array[15777] = 32'hFFFFFFF0;
    // rom_array[15778] = 32'hFFFFFFF0;
    // rom_array[15779] = 32'hFFFFFFF0;
    // rom_array[15780] = 32'hFFFFFFF0;
    // rom_array[15781] = 32'hFFFFFFF1;
    // rom_array[15782] = 32'hFFFFFFF1;
    // rom_array[15783] = 32'hFFFFFFF1;
    // rom_array[15784] = 32'hFFFFFFF1;
    // rom_array[15785] = 32'hFFFFFFF0;
    // rom_array[15786] = 32'hFFFFFFF0;
    // rom_array[15787] = 32'hFFFFFFF0;
    // rom_array[15788] = 32'hFFFFFFF0;
    // rom_array[15789] = 32'hFFFFFFF1;
    // rom_array[15790] = 32'hFFFFFFF1;
    // rom_array[15791] = 32'hFFFFFFF1;
    // rom_array[15792] = 32'hFFFFFFF1;
    // rom_array[15793] = 32'hFFFFFFF0;
    // rom_array[15794] = 32'hFFFFFFF0;
    // rom_array[15795] = 32'hFFFFFFF0;
    // rom_array[15796] = 32'hFFFFFFF0;
    // rom_array[15797] = 32'hFFFFFFF1;
    // rom_array[15798] = 32'hFFFFFFF1;
    // rom_array[15799] = 32'hFFFFFFF1;
    // rom_array[15800] = 32'hFFFFFFF1;
    // rom_array[15801] = 32'hFFFFFFF0;
    // rom_array[15802] = 32'hFFFFFFF0;
    // rom_array[15803] = 32'hFFFFFFF0;
    // rom_array[15804] = 32'hFFFFFFF0;
    // rom_array[15805] = 32'hFFFFFFF1;
    // rom_array[15806] = 32'hFFFFFFF1;
    // rom_array[15807] = 32'hFFFFFFF1;
    // rom_array[15808] = 32'hFFFFFFF1;
    // rom_array[15809] = 32'hFFFFFFF0;
    // rom_array[15810] = 32'hFFFFFFF0;
    // rom_array[15811] = 32'hFFFFFFF0;
    // rom_array[15812] = 32'hFFFFFFF0;
    // rom_array[15813] = 32'hFFFFFFF1;
    // rom_array[15814] = 32'hFFFFFFF1;
    // rom_array[15815] = 32'hFFFFFFF1;
    // rom_array[15816] = 32'hFFFFFFF1;
    // rom_array[15817] = 32'hFFFFFFF1;
    // rom_array[15818] = 32'hFFFFFFF1;
    // rom_array[15819] = 32'hFFFFFFF1;
    // rom_array[15820] = 32'hFFFFFFF1;
    // rom_array[15821] = 32'hFFFFFFF0;
    // rom_array[15822] = 32'hFFFFFFF0;
    // rom_array[15823] = 32'hFFFFFFF0;
    // rom_array[15824] = 32'hFFFFFFF0;
    // rom_array[15825] = 32'hFFFFFFF1;
    // rom_array[15826] = 32'hFFFFFFF1;
    // rom_array[15827] = 32'hFFFFFFF1;
    // rom_array[15828] = 32'hFFFFFFF1;
    // rom_array[15829] = 32'hFFFFFFF0;
    // rom_array[15830] = 32'hFFFFFFF0;
    // rom_array[15831] = 32'hFFFFFFF0;
    // rom_array[15832] = 32'hFFFFFFF0;
    // rom_array[15833] = 32'hFFFFFFF1;
    // rom_array[15834] = 32'hFFFFFFF1;
    // rom_array[15835] = 32'hFFFFFFF1;
    // rom_array[15836] = 32'hFFFFFFF1;
    // rom_array[15837] = 32'hFFFFFFF0;
    // rom_array[15838] = 32'hFFFFFFF0;
    // rom_array[15839] = 32'hFFFFFFF0;
    // rom_array[15840] = 32'hFFFFFFF0;
    // rom_array[15841] = 32'hFFFFFFF1;
    // rom_array[15842] = 32'hFFFFFFF1;
    // rom_array[15843] = 32'hFFFFFFF1;
    // rom_array[15844] = 32'hFFFFFFF1;
    // rom_array[15845] = 32'hFFFFFFF0;
    // rom_array[15846] = 32'hFFFFFFF0;
    // rom_array[15847] = 32'hFFFFFFF0;
    // rom_array[15848] = 32'hFFFFFFF0;
    // rom_array[15849] = 32'hFFFFFFF1;
    // rom_array[15850] = 32'hFFFFFFF1;
    // rom_array[15851] = 32'hFFFFFFF1;
    // rom_array[15852] = 32'hFFFFFFF1;
    // rom_array[15853] = 32'hFFFFFFF0;
    // rom_array[15854] = 32'hFFFFFFF0;
    // rom_array[15855] = 32'hFFFFFFF0;
    // rom_array[15856] = 32'hFFFFFFF0;
    // rom_array[15857] = 32'hFFFFFFF1;
    // rom_array[15858] = 32'hFFFFFFF1;
    // rom_array[15859] = 32'hFFFFFFF1;
    // rom_array[15860] = 32'hFFFFFFF1;
    // rom_array[15861] = 32'hFFFFFFF0;
    // rom_array[15862] = 32'hFFFFFFF0;
    // rom_array[15863] = 32'hFFFFFFF0;
    // rom_array[15864] = 32'hFFFFFFF0;
    // rom_array[15865] = 32'hFFFFFFF1;
    // rom_array[15866] = 32'hFFFFFFF1;
    // rom_array[15867] = 32'hFFFFFFF1;
    // rom_array[15868] = 32'hFFFFFFF1;
    // rom_array[15869] = 32'hFFFFFFF0;
    // rom_array[15870] = 32'hFFFFFFF0;
    // rom_array[15871] = 32'hFFFFFFF0;
    // rom_array[15872] = 32'hFFFFFFF0;
    // rom_array[15873] = 32'hFFFFFFF1;
    // rom_array[15874] = 32'hFFFFFFF1;
    // rom_array[15875] = 32'hFFFFFFF1;
    // rom_array[15876] = 32'hFFFFFFF1;
    // rom_array[15877] = 32'hFFFFFFF0;
    // rom_array[15878] = 32'hFFFFFFF0;
    // rom_array[15879] = 32'hFFFFFFF0;
    // rom_array[15880] = 32'hFFFFFFF0;
    // rom_array[15881] = 32'hFFFFFFF1;
    // rom_array[15882] = 32'hFFFFFFF1;
    // rom_array[15883] = 32'hFFFFFFF1;
    // rom_array[15884] = 32'hFFFFFFF1;
    // rom_array[15885] = 32'hFFFFFFF0;
    // rom_array[15886] = 32'hFFFFFFF0;
    // rom_array[15887] = 32'hFFFFFFF1;
    // rom_array[15888] = 32'hFFFFFFF1;
    // rom_array[15889] = 32'hFFFFFFF1;
    // rom_array[15890] = 32'hFFFFFFF1;
    // rom_array[15891] = 32'hFFFFFFF1;
    // rom_array[15892] = 32'hFFFFFFF1;
    // rom_array[15893] = 32'hFFFFFFF0;
    // rom_array[15894] = 32'hFFFFFFF0;
    // rom_array[15895] = 32'hFFFFFFF1;
    // rom_array[15896] = 32'hFFFFFFF1;
    // rom_array[15897] = 32'hFFFFFFF1;
    // rom_array[15898] = 32'hFFFFFFF1;
    // rom_array[15899] = 32'hFFFFFFF1;
    // rom_array[15900] = 32'hFFFFFFF1;
    // rom_array[15901] = 32'hFFFFFFF1;
    // rom_array[15902] = 32'hFFFFFFF1;
    // rom_array[15903] = 32'hFFFFFFF1;
    // rom_array[15904] = 32'hFFFFFFF1;
    // rom_array[15905] = 32'hFFFFFFF1;
    // rom_array[15906] = 32'hFFFFFFF1;
    // rom_array[15907] = 32'hFFFFFFF1;
    // rom_array[15908] = 32'hFFFFFFF1;
    // rom_array[15909] = 32'hFFFFFFF1;
    // rom_array[15910] = 32'hFFFFFFF1;
    // rom_array[15911] = 32'hFFFFFFF1;
    // rom_array[15912] = 32'hFFFFFFF1;
    // rom_array[15913] = 32'hFFFFFFF0;
    // rom_array[15914] = 32'hFFFFFFF0;
    // rom_array[15915] = 32'hFFFFFFF1;
    // rom_array[15916] = 32'hFFFFFFF1;
    // rom_array[15917] = 32'hFFFFFFF0;
    // rom_array[15918] = 32'hFFFFFFF0;
    // rom_array[15919] = 32'hFFFFFFF1;
    // rom_array[15920] = 32'hFFFFFFF1;
    // rom_array[15921] = 32'hFFFFFFF0;
    // rom_array[15922] = 32'hFFFFFFF0;
    // rom_array[15923] = 32'hFFFFFFF1;
    // rom_array[15924] = 32'hFFFFFFF1;
    // rom_array[15925] = 32'hFFFFFFF0;
    // rom_array[15926] = 32'hFFFFFFF0;
    // rom_array[15927] = 32'hFFFFFFF1;
    // rom_array[15928] = 32'hFFFFFFF1;
    // rom_array[15929] = 32'hFFFFFFF1;
    // rom_array[15930] = 32'hFFFFFFF1;
    // rom_array[15931] = 32'hFFFFFFF1;
    // rom_array[15932] = 32'hFFFFFFF1;
    // rom_array[15933] = 32'hFFFFFFF1;
    // rom_array[15934] = 32'hFFFFFFF1;
    // rom_array[15935] = 32'hFFFFFFF1;
    // rom_array[15936] = 32'hFFFFFFF1;
    // rom_array[15937] = 32'hFFFFFFF1;
    // rom_array[15938] = 32'hFFFFFFF1;
    // rom_array[15939] = 32'hFFFFFFF1;
    // rom_array[15940] = 32'hFFFFFFF1;
    // rom_array[15941] = 32'hFFFFFFF1;
    // rom_array[15942] = 32'hFFFFFFF1;
    // rom_array[15943] = 32'hFFFFFFF1;
    // rom_array[15944] = 32'hFFFFFFF1;
    // rom_array[15945] = 32'hFFFFFFF1;
    // rom_array[15946] = 32'hFFFFFFF1;
    // rom_array[15947] = 32'hFFFFFFF1;
    // rom_array[15948] = 32'hFFFFFFF1;
    // rom_array[15949] = 32'hFFFFFFF1;
    // rom_array[15950] = 32'hFFFFFFF1;
    // rom_array[15951] = 32'hFFFFFFF1;
    // rom_array[15952] = 32'hFFFFFFF1;
    // rom_array[15953] = 32'hFFFFFFF1;
    // rom_array[15954] = 32'hFFFFFFF1;
    // rom_array[15955] = 32'hFFFFFFF1;
    // rom_array[15956] = 32'hFFFFFFF1;
    // rom_array[15957] = 32'hFFFFFFF1;
    // rom_array[15958] = 32'hFFFFFFF1;
    // rom_array[15959] = 32'hFFFFFFF1;
    // rom_array[15960] = 32'hFFFFFFF1;
    // rom_array[15961] = 32'hFFFFFFF0;
    // rom_array[15962] = 32'hFFFFFFF0;
    // rom_array[15963] = 32'hFFFFFFF1;
    // rom_array[15964] = 32'hFFFFFFF1;
    // rom_array[15965] = 32'hFFFFFFF0;
    // rom_array[15966] = 32'hFFFFFFF0;
    // rom_array[15967] = 32'hFFFFFFF1;
    // rom_array[15968] = 32'hFFFFFFF1;
    // rom_array[15969] = 32'hFFFFFFF0;
    // rom_array[15970] = 32'hFFFFFFF0;
    // rom_array[15971] = 32'hFFFFFFF1;
    // rom_array[15972] = 32'hFFFFFFF1;
    // rom_array[15973] = 32'hFFFFFFF0;
    // rom_array[15974] = 32'hFFFFFFF0;
    // rom_array[15975] = 32'hFFFFFFF1;
    // rom_array[15976] = 32'hFFFFFFF1;
    // rom_array[15977] = 32'hFFFFFFF0;
    // rom_array[15978] = 32'hFFFFFFF0;
    // rom_array[15979] = 32'hFFFFFFF1;
    // rom_array[15980] = 32'hFFFFFFF1;
    // rom_array[15981] = 32'hFFFFFFF0;
    // rom_array[15982] = 32'hFFFFFFF0;
    // rom_array[15983] = 32'hFFFFFFF1;
    // rom_array[15984] = 32'hFFFFFFF1;
    // rom_array[15985] = 32'hFFFFFFF0;
    // rom_array[15986] = 32'hFFFFFFF0;
    // rom_array[15987] = 32'hFFFFFFF1;
    // rom_array[15988] = 32'hFFFFFFF1;
    // rom_array[15989] = 32'hFFFFFFF0;
    // rom_array[15990] = 32'hFFFFFFF0;
    // rom_array[15991] = 32'hFFFFFFF1;
    // rom_array[15992] = 32'hFFFFFFF1;
    // rom_array[15993] = 32'hFFFFFFF0;
    // rom_array[15994] = 32'hFFFFFFF0;
    // rom_array[15995] = 32'hFFFFFFF1;
    // rom_array[15996] = 32'hFFFFFFF1;
    // rom_array[15997] = 32'hFFFFFFF0;
    // rom_array[15998] = 32'hFFFFFFF0;
    // rom_array[15999] = 32'hFFFFFFF1;
    // rom_array[16000] = 32'hFFFFFFF1;
    // rom_array[16001] = 32'hFFFFFFF0;
    // rom_array[16002] = 32'hFFFFFFF0;
    // rom_array[16003] = 32'hFFFFFFF1;
    // rom_array[16004] = 32'hFFFFFFF1;
    // rom_array[16005] = 32'hFFFFFFF0;
    // rom_array[16006] = 32'hFFFFFFF0;
    // rom_array[16007] = 32'hFFFFFFF1;
    // rom_array[16008] = 32'hFFFFFFF1;
    // rom_array[16009] = 32'hFFFFFFF0;
    // rom_array[16010] = 32'hFFFFFFF0;
    // rom_array[16011] = 32'hFFFFFFF1;
    // rom_array[16012] = 32'hFFFFFFF1;
    // rom_array[16013] = 32'hFFFFFFF0;
    // rom_array[16014] = 32'hFFFFFFF0;
    // rom_array[16015] = 32'hFFFFFFF1;
    // rom_array[16016] = 32'hFFFFFFF1;
    // rom_array[16017] = 32'hFFFFFFF0;
    // rom_array[16018] = 32'hFFFFFFF0;
    // rom_array[16019] = 32'hFFFFFFF1;
    // rom_array[16020] = 32'hFFFFFFF1;
    // rom_array[16021] = 32'hFFFFFFF0;
    // rom_array[16022] = 32'hFFFFFFF0;
    // rom_array[16023] = 32'hFFFFFFF1;
    // rom_array[16024] = 32'hFFFFFFF1;
    // rom_array[16025] = 32'hFFFFFFF0;
    // rom_array[16026] = 32'hFFFFFFF0;
    // rom_array[16027] = 32'hFFFFFFF1;
    // rom_array[16028] = 32'hFFFFFFF1;
    // rom_array[16029] = 32'hFFFFFFF0;
    // rom_array[16030] = 32'hFFFFFFF0;
    // rom_array[16031] = 32'hFFFFFFF1;
    // rom_array[16032] = 32'hFFFFFFF1;
    // rom_array[16033] = 32'hFFFFFFF0;
    // rom_array[16034] = 32'hFFFFFFF0;
    // rom_array[16035] = 32'hFFFFFFF1;
    // rom_array[16036] = 32'hFFFFFFF1;
    // rom_array[16037] = 32'hFFFFFFF0;
    // rom_array[16038] = 32'hFFFFFFF0;
    // rom_array[16039] = 32'hFFFFFFF1;
    // rom_array[16040] = 32'hFFFFFFF1;
    // rom_array[16041] = 32'hFFFFFFF0;
    // rom_array[16042] = 32'hFFFFFFF0;
    // rom_array[16043] = 32'hFFFFFFF1;
    // rom_array[16044] = 32'hFFFFFFF1;
    // rom_array[16045] = 32'hFFFFFFF0;
    // rom_array[16046] = 32'hFFFFFFF0;
    // rom_array[16047] = 32'hFFFFFFF1;
    // rom_array[16048] = 32'hFFFFFFF1;
    // rom_array[16049] = 32'hFFFFFFF0;
    // rom_array[16050] = 32'hFFFFFFF0;
    // rom_array[16051] = 32'hFFFFFFF1;
    // rom_array[16052] = 32'hFFFFFFF1;
    // rom_array[16053] = 32'hFFFFFFF0;
    // rom_array[16054] = 32'hFFFFFFF0;
    // rom_array[16055] = 32'hFFFFFFF1;
    // rom_array[16056] = 32'hFFFFFFF1;
    // rom_array[16057] = 32'hFFFFFFF0;
    // rom_array[16058] = 32'hFFFFFFF0;
    // rom_array[16059] = 32'hFFFFFFF0;
    // rom_array[16060] = 32'hFFFFFFF0;
    // rom_array[16061] = 32'hFFFFFFF0;
    // rom_array[16062] = 32'hFFFFFFF0;
    // rom_array[16063] = 32'hFFFFFFF1;
    // rom_array[16064] = 32'hFFFFFFF1;
    // rom_array[16065] = 32'hFFFFFFF0;
    // rom_array[16066] = 32'hFFFFFFF0;
    // rom_array[16067] = 32'hFFFFFFF0;
    // rom_array[16068] = 32'hFFFFFFF0;
    // rom_array[16069] = 32'hFFFFFFF0;
    // rom_array[16070] = 32'hFFFFFFF0;
    // rom_array[16071] = 32'hFFFFFFF1;
    // rom_array[16072] = 32'hFFFFFFF1;
    // rom_array[16073] = 32'hFFFFFFF0;
    // rom_array[16074] = 32'hFFFFFFF0;
    // rom_array[16075] = 32'hFFFFFFF1;
    // rom_array[16076] = 32'hFFFFFFF1;
    // rom_array[16077] = 32'hFFFFFFF0;
    // rom_array[16078] = 32'hFFFFFFF0;
    // rom_array[16079] = 32'hFFFFFFF0;
    // rom_array[16080] = 32'hFFFFFFF0;
    // rom_array[16081] = 32'hFFFFFFF0;
    // rom_array[16082] = 32'hFFFFFFF0;
    // rom_array[16083] = 32'hFFFFFFF1;
    // rom_array[16084] = 32'hFFFFFFF1;
    // rom_array[16085] = 32'hFFFFFFF0;
    // rom_array[16086] = 32'hFFFFFFF0;
    // rom_array[16087] = 32'hFFFFFFF0;
    // rom_array[16088] = 32'hFFFFFFF0;
    // rom_array[16089] = 32'hFFFFFFF1;
    // rom_array[16090] = 32'hFFFFFFF1;
    // rom_array[16091] = 32'hFFFFFFF1;
    // rom_array[16092] = 32'hFFFFFFF1;
    // rom_array[16093] = 32'hFFFFFFF0;
    // rom_array[16094] = 32'hFFFFFFF0;
    // rom_array[16095] = 32'hFFFFFFF0;
    // rom_array[16096] = 32'hFFFFFFF0;
    // rom_array[16097] = 32'hFFFFFFF1;
    // rom_array[16098] = 32'hFFFFFFF1;
    // rom_array[16099] = 32'hFFFFFFF1;
    // rom_array[16100] = 32'hFFFFFFF1;
    // rom_array[16101] = 32'hFFFFFFF0;
    // rom_array[16102] = 32'hFFFFFFF0;
    // rom_array[16103] = 32'hFFFFFFF0;
    // rom_array[16104] = 32'hFFFFFFF0;
    // rom_array[16105] = 32'hFFFFFFF1;
    // rom_array[16106] = 32'hFFFFFFF1;
    // rom_array[16107] = 32'hFFFFFFF1;
    // rom_array[16108] = 32'hFFFFFFF1;
    // rom_array[16109] = 32'hFFFFFFF0;
    // rom_array[16110] = 32'hFFFFFFF0;
    // rom_array[16111] = 32'hFFFFFFF0;
    // rom_array[16112] = 32'hFFFFFFF0;
    // rom_array[16113] = 32'hFFFFFFF1;
    // rom_array[16114] = 32'hFFFFFFF1;
    // rom_array[16115] = 32'hFFFFFFF1;
    // rom_array[16116] = 32'hFFFFFFF1;
    // rom_array[16117] = 32'hFFFFFFF0;
    // rom_array[16118] = 32'hFFFFFFF0;
    // rom_array[16119] = 32'hFFFFFFF0;
    // rom_array[16120] = 32'hFFFFFFF0;
    // rom_array[16121] = 32'hFFFFFFF1;
    // rom_array[16122] = 32'hFFFFFFF1;
    // rom_array[16123] = 32'hFFFFFFF1;
    // rom_array[16124] = 32'hFFFFFFF1;
    // rom_array[16125] = 32'hFFFFFFF0;
    // rom_array[16126] = 32'hFFFFFFF0;
    // rom_array[16127] = 32'hFFFFFFF1;
    // rom_array[16128] = 32'hFFFFFFF1;
    // rom_array[16129] = 32'hFFFFFFF1;
    // rom_array[16130] = 32'hFFFFFFF1;
    // rom_array[16131] = 32'hFFFFFFF1;
    // rom_array[16132] = 32'hFFFFFFF1;
    // rom_array[16133] = 32'hFFFFFFF0;
    // rom_array[16134] = 32'hFFFFFFF0;
    // rom_array[16135] = 32'hFFFFFFF1;
    // rom_array[16136] = 32'hFFFFFFF1;
    // rom_array[16137] = 32'hFFFFFFF0;
    // rom_array[16138] = 32'hFFFFFFF0;
    // rom_array[16139] = 32'hFFFFFFF1;
    // rom_array[16140] = 32'hFFFFFFF1;
    // rom_array[16141] = 32'hFFFFFFF0;
    // rom_array[16142] = 32'hFFFFFFF0;
    // rom_array[16143] = 32'hFFFFFFF1;
    // rom_array[16144] = 32'hFFFFFFF1;
    // rom_array[16145] = 32'hFFFFFFF0;
    // rom_array[16146] = 32'hFFFFFFF0;
    // rom_array[16147] = 32'hFFFFFFF1;
    // rom_array[16148] = 32'hFFFFFFF1;
    // rom_array[16149] = 32'hFFFFFFF0;
    // rom_array[16150] = 32'hFFFFFFF0;
    // rom_array[16151] = 32'hFFFFFFF1;
    // rom_array[16152] = 32'hFFFFFFF1;
    // rom_array[16153] = 32'hFFFFFFF0;
    // rom_array[16154] = 32'hFFFFFFF0;
    // rom_array[16155] = 32'hFFFFFFF1;
    // rom_array[16156] = 32'hFFFFFFF1;
    // rom_array[16157] = 32'hFFFFFFF0;
    // rom_array[16158] = 32'hFFFFFFF0;
    // rom_array[16159] = 32'hFFFFFFF1;
    // rom_array[16160] = 32'hFFFFFFF1;
    // rom_array[16161] = 32'hFFFFFFF0;
    // rom_array[16162] = 32'hFFFFFFF0;
    // rom_array[16163] = 32'hFFFFFFF1;
    // rom_array[16164] = 32'hFFFFFFF1;
    // rom_array[16165] = 32'hFFFFFFF0;
    // rom_array[16166] = 32'hFFFFFFF0;
    // rom_array[16167] = 32'hFFFFFFF1;
    // rom_array[16168] = 32'hFFFFFFF1;
    // rom_array[16169] = 32'hFFFFFFF0;
    // rom_array[16170] = 32'hFFFFFFF0;
    // rom_array[16171] = 32'hFFFFFFF1;
    // rom_array[16172] = 32'hFFFFFFF1;
    // rom_array[16173] = 32'hFFFFFFF0;
    // rom_array[16174] = 32'hFFFFFFF0;
    // rom_array[16175] = 32'hFFFFFFF0;
    // rom_array[16176] = 32'hFFFFFFF0;
    // rom_array[16177] = 32'hFFFFFFF0;
    // rom_array[16178] = 32'hFFFFFFF0;
    // rom_array[16179] = 32'hFFFFFFF1;
    // rom_array[16180] = 32'hFFFFFFF1;
    // rom_array[16181] = 32'hFFFFFFF0;
    // rom_array[16182] = 32'hFFFFFFF0;
    // rom_array[16183] = 32'hFFFFFFF0;
    // rom_array[16184] = 32'hFFFFFFF0;
    // rom_array[16185] = 32'hFFFFFFF0;
    // rom_array[16186] = 32'hFFFFFFF0;
    // rom_array[16187] = 32'hFFFFFFF0;
    // rom_array[16188] = 32'hFFFFFFF0;
    // rom_array[16189] = 32'hFFFFFFF0;
    // rom_array[16190] = 32'hFFFFFFF0;
    // rom_array[16191] = 32'hFFFFFFF1;
    // rom_array[16192] = 32'hFFFFFFF1;
    // rom_array[16193] = 32'hFFFFFFF0;
    // rom_array[16194] = 32'hFFFFFFF0;
    // rom_array[16195] = 32'hFFFFFFF0;
    // rom_array[16196] = 32'hFFFFFFF0;
    // rom_array[16197] = 32'hFFFFFFF0;
    // rom_array[16198] = 32'hFFFFFFF0;
    // rom_array[16199] = 32'hFFFFFFF1;
    // rom_array[16200] = 32'hFFFFFFF1;
    // rom_array[16201] = 32'hFFFFFFF0;
    // rom_array[16202] = 32'hFFFFFFF0;
    // rom_array[16203] = 32'hFFFFFFF0;
    // rom_array[16204] = 32'hFFFFFFF0;
    // rom_array[16205] = 32'hFFFFFFF1;
    // rom_array[16206] = 32'hFFFFFFF1;
    // rom_array[16207] = 32'hFFFFFFF1;
    // rom_array[16208] = 32'hFFFFFFF1;
    // rom_array[16209] = 32'hFFFFFFF0;
    // rom_array[16210] = 32'hFFFFFFF0;
    // rom_array[16211] = 32'hFFFFFFF0;
    // rom_array[16212] = 32'hFFFFFFF0;
    // rom_array[16213] = 32'hFFFFFFF1;
    // rom_array[16214] = 32'hFFFFFFF1;
    // rom_array[16215] = 32'hFFFFFFF1;
    // rom_array[16216] = 32'hFFFFFFF1;
    // rom_array[16217] = 32'hFFFFFFF0;
    // rom_array[16218] = 32'hFFFFFFF0;
    // rom_array[16219] = 32'hFFFFFFF1;
    // rom_array[16220] = 32'hFFFFFFF1;
    // rom_array[16221] = 32'hFFFFFFF0;
    // rom_array[16222] = 32'hFFFFFFF0;
    // rom_array[16223] = 32'hFFFFFFF1;
    // rom_array[16224] = 32'hFFFFFFF1;
    // rom_array[16225] = 32'hFFFFFFF0;
    // rom_array[16226] = 32'hFFFFFFF0;
    // rom_array[16227] = 32'hFFFFFFF1;
    // rom_array[16228] = 32'hFFFFFFF1;
    // rom_array[16229] = 32'hFFFFFFF0;
    // rom_array[16230] = 32'hFFFFFFF0;
    // rom_array[16231] = 32'hFFFFFFF1;
    // rom_array[16232] = 32'hFFFFFFF1;
    // rom_array[16233] = 32'hFFFFFFF0;
    // rom_array[16234] = 32'hFFFFFFF0;
    // rom_array[16235] = 32'hFFFFFFF0;
    // rom_array[16236] = 32'hFFFFFFF0;
    // rom_array[16237] = 32'hFFFFFFF1;
    // rom_array[16238] = 32'hFFFFFFF1;
    // rom_array[16239] = 32'hFFFFFFF1;
    // rom_array[16240] = 32'hFFFFFFF1;
    // rom_array[16241] = 32'hFFFFFFF0;
    // rom_array[16242] = 32'hFFFFFFF0;
    // rom_array[16243] = 32'hFFFFFFF0;
    // rom_array[16244] = 32'hFFFFFFF0;
    // rom_array[16245] = 32'hFFFFFFF1;
    // rom_array[16246] = 32'hFFFFFFF1;
    // rom_array[16247] = 32'hFFFFFFF1;
    // rom_array[16248] = 32'hFFFFFFF1;
    // rom_array[16249] = 32'hFFFFFFF0;
    // rom_array[16250] = 32'hFFFFFFF0;
    // rom_array[16251] = 32'hFFFFFFF0;
    // rom_array[16252] = 32'hFFFFFFF0;
    // rom_array[16253] = 32'hFFFFFFF1;
    // rom_array[16254] = 32'hFFFFFFF1;
    // rom_array[16255] = 32'hFFFFFFF1;
    // rom_array[16256] = 32'hFFFFFFF1;
    // rom_array[16257] = 32'hFFFFFFF0;
    // rom_array[16258] = 32'hFFFFFFF0;
    // rom_array[16259] = 32'hFFFFFFF0;
    // rom_array[16260] = 32'hFFFFFFF0;
    // rom_array[16261] = 32'hFFFFFFF1;
    // rom_array[16262] = 32'hFFFFFFF1;
    // rom_array[16263] = 32'hFFFFFFF1;
    // rom_array[16264] = 32'hFFFFFFF1;
    // rom_array[16265] = 32'hFFFFFFF0;
    // rom_array[16266] = 32'hFFFFFFF0;
    // rom_array[16267] = 32'hFFFFFFF1;
    // rom_array[16268] = 32'hFFFFFFF1;
    // rom_array[16269] = 32'hFFFFFFF0;
    // rom_array[16270] = 32'hFFFFFFF0;
    // rom_array[16271] = 32'hFFFFFFF1;
    // rom_array[16272] = 32'hFFFFFFF1;
    // rom_array[16273] = 32'hFFFFFFF0;
    // rom_array[16274] = 32'hFFFFFFF0;
    // rom_array[16275] = 32'hFFFFFFF1;
    // rom_array[16276] = 32'hFFFFFFF1;
    // rom_array[16277] = 32'hFFFFFFF0;
    // rom_array[16278] = 32'hFFFFFFF0;
    // rom_array[16279] = 32'hFFFFFFF1;
    // rom_array[16280] = 32'hFFFFFFF1;
    // rom_array[16281] = 32'hFFFFFFF0;
    // rom_array[16282] = 32'hFFFFFFF0;
    // rom_array[16283] = 32'hFFFFFFF1;
    // rom_array[16284] = 32'hFFFFFFF1;
    // rom_array[16285] = 32'hFFFFFFF0;
    // rom_array[16286] = 32'hFFFFFFF0;
    // rom_array[16287] = 32'hFFFFFFF1;
    // rom_array[16288] = 32'hFFFFFFF1;
    // rom_array[16289] = 32'hFFFFFFF0;
    // rom_array[16290] = 32'hFFFFFFF0;
    // rom_array[16291] = 32'hFFFFFFF1;
    // rom_array[16292] = 32'hFFFFFFF1;
    // rom_array[16293] = 32'hFFFFFFF0;
    // rom_array[16294] = 32'hFFFFFFF0;
    // rom_array[16295] = 32'hFFFFFFF1;
    // rom_array[16296] = 32'hFFFFFFF1;
    // rom_array[16297] = 32'hFFFFFFF0;
    // rom_array[16298] = 32'hFFFFFFF0;
    // rom_array[16299] = 32'hFFFFFFF1;
    // rom_array[16300] = 32'hFFFFFFF1;
    // rom_array[16301] = 32'hFFFFFFF0;
    // rom_array[16302] = 32'hFFFFFFF0;
    // rom_array[16303] = 32'hFFFFFFF1;
    // rom_array[16304] = 32'hFFFFFFF1;
    // rom_array[16305] = 32'hFFFFFFF0;
    // rom_array[16306] = 32'hFFFFFFF0;
    // rom_array[16307] = 32'hFFFFFFF1;
    // rom_array[16308] = 32'hFFFFFFF1;
    // rom_array[16309] = 32'hFFFFFFF0;
    // rom_array[16310] = 32'hFFFFFFF0;
    // rom_array[16311] = 32'hFFFFFFF1;
    // rom_array[16312] = 32'hFFFFFFF1;
    // rom_array[16313] = 32'hFFFFFFF1;
    // rom_array[16314] = 32'hFFFFFFF1;
    // rom_array[16315] = 32'hFFFFFFF1;
    // rom_array[16316] = 32'hFFFFFFF1;
    // rom_array[16317] = 32'hFFFFFFF1;
    // rom_array[16318] = 32'hFFFFFFF1;
    // rom_array[16319] = 32'hFFFFFFF1;
    // rom_array[16320] = 32'hFFFFFFF1;
    // rom_array[16321] = 32'hFFFFFFF1;
    // rom_array[16322] = 32'hFFFFFFF1;
    // rom_array[16323] = 32'hFFFFFFF1;
    // rom_array[16324] = 32'hFFFFFFF1;
    // rom_array[16325] = 32'hFFFFFFF1;
    // rom_array[16326] = 32'hFFFFFFF1;
    // rom_array[16327] = 32'hFFFFFFF1;
    // rom_array[16328] = 32'hFFFFFFF1;
    // rom_array[16329] = 32'hFFFFFFF0;
    // rom_array[16330] = 32'hFFFFFFF0;
    // rom_array[16331] = 32'hFFFFFFF1;
    // rom_array[16332] = 32'hFFFFFFF1;
    // rom_array[16333] = 32'hFFFFFFF0;
    // rom_array[16334] = 32'hFFFFFFF0;
    // rom_array[16335] = 32'hFFFFFFF1;
    // rom_array[16336] = 32'hFFFFFFF1;
    // rom_array[16337] = 32'hFFFFFFF0;
    // rom_array[16338] = 32'hFFFFFFF0;
    // rom_array[16339] = 32'hFFFFFFF1;
    // rom_array[16340] = 32'hFFFFFFF1;
    // rom_array[16341] = 32'hFFFFFFF0;
    // rom_array[16342] = 32'hFFFFFFF0;
    // rom_array[16343] = 32'hFFFFFFF1;
    // rom_array[16344] = 32'hFFFFFFF1;
    // rom_array[16345] = 32'hFFFFFFF1;
    // rom_array[16346] = 32'hFFFFFFF1;
    // rom_array[16347] = 32'hFFFFFFF1;
    // rom_array[16348] = 32'hFFFFFFF1;
    // rom_array[16349] = 32'hFFFFFFF1;
    // rom_array[16350] = 32'hFFFFFFF1;
    // rom_array[16351] = 32'hFFFFFFF1;
    // rom_array[16352] = 32'hFFFFFFF1;
    // rom_array[16353] = 32'hFFFFFFF1;
    // rom_array[16354] = 32'hFFFFFFF1;
    // rom_array[16355] = 32'hFFFFFFF1;
    // rom_array[16356] = 32'hFFFFFFF1;
    // rom_array[16357] = 32'hFFFFFFF1;
    // rom_array[16358] = 32'hFFFFFFF1;
    // rom_array[16359] = 32'hFFFFFFF1;
    // rom_array[16360] = 32'hFFFFFFF1;
    // rom_array[16361] = 32'hFFFFFFF1;
    // rom_array[16362] = 32'hFFFFFFF1;
    // rom_array[16363] = 32'hFFFFFFF1;
    // rom_array[16364] = 32'hFFFFFFF1;
    // rom_array[16365] = 32'hFFFFFFF1;
    // rom_array[16366] = 32'hFFFFFFF1;
    // rom_array[16367] = 32'hFFFFFFF1;
    // rom_array[16368] = 32'hFFFFFFF1;
    // rom_array[16369] = 32'hFFFFFFF1;
    // rom_array[16370] = 32'hFFFFFFF1;
    // rom_array[16371] = 32'hFFFFFFF1;
    // rom_array[16372] = 32'hFFFFFFF1;
    // rom_array[16373] = 32'hFFFFFFF1;
    // rom_array[16374] = 32'hFFFFFFF1;
    // rom_array[16375] = 32'hFFFFFFF1;
    // rom_array[16376] = 32'hFFFFFFF1;
    // rom_array[16377] = 32'hFFFFFFF0;
    // rom_array[16378] = 32'hFFFFFFF0;
    // rom_array[16379] = 32'hFFFFFFF0;
    // rom_array[16380] = 32'hFFFFFFF0;
    // rom_array[16381] = 32'hFFFFFFF1;
    // rom_array[16382] = 32'hFFFFFFF1;
    // rom_array[16383] = 32'hFFFFFFF1;
    // rom_array[16384] = 32'hFFFFFFF1;
    // rom_array[16385] = 32'hFFFFFFF0;
    // rom_array[16386] = 32'hFFFFFFF0;
    // rom_array[16387] = 32'hFFFFFFF0;
    // rom_array[16388] = 32'hFFFFFFF0;
    // rom_array[16389] = 32'hFFFFFFF1;
    // rom_array[16390] = 32'hFFFFFFF1;
    // rom_array[16391] = 32'hFFFFFFF1;
    // rom_array[16392] = 32'hFFFFFFF1;
    // rom_array[16393] = 32'hFFFFFFF0;
    // rom_array[16394] = 32'hFFFFFFF0;
    // rom_array[16395] = 32'hFFFFFFF0;
    // rom_array[16396] = 32'hFFFFFFF0;
    // rom_array[16397] = 32'hFFFFFFF1;
    // rom_array[16398] = 32'hFFFFFFF1;
    // rom_array[16399] = 32'hFFFFFFF1;
    // rom_array[16400] = 32'hFFFFFFF1;
    // rom_array[16401] = 32'hFFFFFFF0;
    // rom_array[16402] = 32'hFFFFFFF0;
    // rom_array[16403] = 32'hFFFFFFF0;
    // rom_array[16404] = 32'hFFFFFFF0;
    // rom_array[16405] = 32'hFFFFFFF1;
    // rom_array[16406] = 32'hFFFFFFF1;
    // rom_array[16407] = 32'hFFFFFFF1;
    // rom_array[16408] = 32'hFFFFFFF1;
    // rom_array[16409] = 32'hFFFFFFF0;
    // rom_array[16410] = 32'hFFFFFFF0;
    // rom_array[16411] = 32'hFFFFFFF0;
    // rom_array[16412] = 32'hFFFFFFF0;
    // rom_array[16413] = 32'hFFFFFFF1;
    // rom_array[16414] = 32'hFFFFFFF1;
    // rom_array[16415] = 32'hFFFFFFF1;
    // rom_array[16416] = 32'hFFFFFFF1;
    // rom_array[16417] = 32'hFFFFFFF0;
    // rom_array[16418] = 32'hFFFFFFF0;
    // rom_array[16419] = 32'hFFFFFFF0;
    // rom_array[16420] = 32'hFFFFFFF0;
    // rom_array[16421] = 32'hFFFFFFF1;
    // rom_array[16422] = 32'hFFFFFFF1;
    // rom_array[16423] = 32'hFFFFFFF1;
    // rom_array[16424] = 32'hFFFFFFF1;
    // rom_array[16425] = 32'hFFFFFFF0;
    // rom_array[16426] = 32'hFFFFFFF0;
    // rom_array[16427] = 32'hFFFFFFF0;
    // rom_array[16428] = 32'hFFFFFFF0;
    // rom_array[16429] = 32'hFFFFFFF1;
    // rom_array[16430] = 32'hFFFFFFF1;
    // rom_array[16431] = 32'hFFFFFFF1;
    // rom_array[16432] = 32'hFFFFFFF1;
    // rom_array[16433] = 32'hFFFFFFF0;
    // rom_array[16434] = 32'hFFFFFFF0;
    // rom_array[16435] = 32'hFFFFFFF0;
    // rom_array[16436] = 32'hFFFFFFF0;
    // rom_array[16437] = 32'hFFFFFFF1;
    // rom_array[16438] = 32'hFFFFFFF1;
    // rom_array[16439] = 32'hFFFFFFF1;
    // rom_array[16440] = 32'hFFFFFFF1;
    // rom_array[16441] = 32'hFFFFFFF0;
    // rom_array[16442] = 32'hFFFFFFF0;
    // rom_array[16443] = 32'hFFFFFFF0;
    // rom_array[16444] = 32'hFFFFFFF0;
    // rom_array[16445] = 32'hFFFFFFF1;
    // rom_array[16446] = 32'hFFFFFFF1;
    // rom_array[16447] = 32'hFFFFFFF1;
    // rom_array[16448] = 32'hFFFFFFF1;
    // rom_array[16449] = 32'hFFFFFFF0;
    // rom_array[16450] = 32'hFFFFFFF0;
    // rom_array[16451] = 32'hFFFFFFF0;
    // rom_array[16452] = 32'hFFFFFFF0;
    // rom_array[16453] = 32'hFFFFFFF1;
    // rom_array[16454] = 32'hFFFFFFF1;
    // rom_array[16455] = 32'hFFFFFFF1;
    // rom_array[16456] = 32'hFFFFFFF1;
    // rom_array[16457] = 32'hFFFFFFF0;
    // rom_array[16458] = 32'hFFFFFFF0;
    // rom_array[16459] = 32'hFFFFFFF0;
    // rom_array[16460] = 32'hFFFFFFF0;
    // rom_array[16461] = 32'hFFFFFFF1;
    // rom_array[16462] = 32'hFFFFFFF1;
    // rom_array[16463] = 32'hFFFFFFF1;
    // rom_array[16464] = 32'hFFFFFFF1;
    // rom_array[16465] = 32'hFFFFFFF0;
    // rom_array[16466] = 32'hFFFFFFF0;
    // rom_array[16467] = 32'hFFFFFFF0;
    // rom_array[16468] = 32'hFFFFFFF0;
    // rom_array[16469] = 32'hFFFFFFF1;
    // rom_array[16470] = 32'hFFFFFFF1;
    // rom_array[16471] = 32'hFFFFFFF1;
    // rom_array[16472] = 32'hFFFFFFF1;
    // rom_array[16473] = 32'hFFFFFFF0;
    // rom_array[16474] = 32'hFFFFFFF0;
    // rom_array[16475] = 32'hFFFFFFF0;
    // rom_array[16476] = 32'hFFFFFFF0;
    // rom_array[16477] = 32'hFFFFFFF1;
    // rom_array[16478] = 32'hFFFFFFF1;
    // rom_array[16479] = 32'hFFFFFFF1;
    // rom_array[16480] = 32'hFFFFFFF1;
    // rom_array[16481] = 32'hFFFFFFF0;
    // rom_array[16482] = 32'hFFFFFFF0;
    // rom_array[16483] = 32'hFFFFFFF0;
    // rom_array[16484] = 32'hFFFFFFF0;
    // rom_array[16485] = 32'hFFFFFFF1;
    // rom_array[16486] = 32'hFFFFFFF1;
    // rom_array[16487] = 32'hFFFFFFF1;
    // rom_array[16488] = 32'hFFFFFFF1;
    // rom_array[16489] = 32'hFFFFFFF0;
    // rom_array[16490] = 32'hFFFFFFF0;
    // rom_array[16491] = 32'hFFFFFFF0;
    // rom_array[16492] = 32'hFFFFFFF0;
    // rom_array[16493] = 32'hFFFFFFF1;
    // rom_array[16494] = 32'hFFFFFFF1;
    // rom_array[16495] = 32'hFFFFFFF1;
    // rom_array[16496] = 32'hFFFFFFF1;
    // rom_array[16497] = 32'hFFFFFFF0;
    // rom_array[16498] = 32'hFFFFFFF0;
    // rom_array[16499] = 32'hFFFFFFF0;
    // rom_array[16500] = 32'hFFFFFFF0;
    // rom_array[16501] = 32'hFFFFFFF1;
    // rom_array[16502] = 32'hFFFFFFF1;
    // rom_array[16503] = 32'hFFFFFFF1;
    // rom_array[16504] = 32'hFFFFFFF1;
    // rom_array[16505] = 32'hFFFFFFF1;
    // rom_array[16506] = 32'hFFFFFFF1;
    // rom_array[16507] = 32'hFFFFFFF1;
    // rom_array[16508] = 32'hFFFFFFF1;
    // rom_array[16509] = 32'hFFFFFFF1;
    // rom_array[16510] = 32'hFFFFFFF1;
    // rom_array[16511] = 32'hFFFFFFF1;
    // rom_array[16512] = 32'hFFFFFFF1;
    // rom_array[16513] = 32'hFFFFFFF1;
    // rom_array[16514] = 32'hFFFFFFF1;
    // rom_array[16515] = 32'hFFFFFFF1;
    // rom_array[16516] = 32'hFFFFFFF1;
    // rom_array[16517] = 32'hFFFFFFF1;
    // rom_array[16518] = 32'hFFFFFFF1;
    // rom_array[16519] = 32'hFFFFFFF1;
    // rom_array[16520] = 32'hFFFFFFF1;
    // rom_array[16521] = 32'hFFFFFFF1;
    // rom_array[16522] = 32'hFFFFFFF1;
    // rom_array[16523] = 32'hFFFFFFF1;
    // rom_array[16524] = 32'hFFFFFFF1;
    // rom_array[16525] = 32'hFFFFFFF0;
    // rom_array[16526] = 32'hFFFFFFF0;
    // rom_array[16527] = 32'hFFFFFFF0;
    // rom_array[16528] = 32'hFFFFFFF0;
    // rom_array[16529] = 32'hFFFFFFF1;
    // rom_array[16530] = 32'hFFFFFFF1;
    // rom_array[16531] = 32'hFFFFFFF1;
    // rom_array[16532] = 32'hFFFFFFF1;
    // rom_array[16533] = 32'hFFFFFFF0;
    // rom_array[16534] = 32'hFFFFFFF0;
    // rom_array[16535] = 32'hFFFFFFF0;
    // rom_array[16536] = 32'hFFFFFFF0;
    // rom_array[16537] = 32'hFFFFFFF1;
    // rom_array[16538] = 32'hFFFFFFF1;
    // rom_array[16539] = 32'hFFFFFFF1;
    // rom_array[16540] = 32'hFFFFFFF1;
    // rom_array[16541] = 32'hFFFFFFF1;
    // rom_array[16542] = 32'hFFFFFFF1;
    // rom_array[16543] = 32'hFFFFFFF1;
    // rom_array[16544] = 32'hFFFFFFF1;
    // rom_array[16545] = 32'hFFFFFFF1;
    // rom_array[16546] = 32'hFFFFFFF1;
    // rom_array[16547] = 32'hFFFFFFF1;
    // rom_array[16548] = 32'hFFFFFFF1;
    // rom_array[16549] = 32'hFFFFFFF1;
    // rom_array[16550] = 32'hFFFFFFF1;
    // rom_array[16551] = 32'hFFFFFFF1;
    // rom_array[16552] = 32'hFFFFFFF1;
    // rom_array[16553] = 32'hFFFFFFF1;
    // rom_array[16554] = 32'hFFFFFFF1;
    // rom_array[16555] = 32'hFFFFFFF1;
    // rom_array[16556] = 32'hFFFFFFF1;
    // rom_array[16557] = 32'hFFFFFFF0;
    // rom_array[16558] = 32'hFFFFFFF0;
    // rom_array[16559] = 32'hFFFFFFF0;
    // rom_array[16560] = 32'hFFFFFFF0;
    // rom_array[16561] = 32'hFFFFFFF1;
    // rom_array[16562] = 32'hFFFFFFF1;
    // rom_array[16563] = 32'hFFFFFFF1;
    // rom_array[16564] = 32'hFFFFFFF1;
    // rom_array[16565] = 32'hFFFFFFF0;
    // rom_array[16566] = 32'hFFFFFFF0;
    // rom_array[16567] = 32'hFFFFFFF0;
    // rom_array[16568] = 32'hFFFFFFF0;
    // rom_array[16569] = 32'hFFFFFFF1;
    // rom_array[16570] = 32'hFFFFFFF1;
    // rom_array[16571] = 32'hFFFFFFF1;
    // rom_array[16572] = 32'hFFFFFFF1;
    // rom_array[16573] = 32'hFFFFFFF0;
    // rom_array[16574] = 32'hFFFFFFF0;
    // rom_array[16575] = 32'hFFFFFFF0;
    // rom_array[16576] = 32'hFFFFFFF0;
    // rom_array[16577] = 32'hFFFFFFF1;
    // rom_array[16578] = 32'hFFFFFFF1;
    // rom_array[16579] = 32'hFFFFFFF1;
    // rom_array[16580] = 32'hFFFFFFF1;
    // rom_array[16581] = 32'hFFFFFFF0;
    // rom_array[16582] = 32'hFFFFFFF0;
    // rom_array[16583] = 32'hFFFFFFF0;
    // rom_array[16584] = 32'hFFFFFFF0;
    // rom_array[16585] = 32'hFFFFFFF1;
    // rom_array[16586] = 32'hFFFFFFF1;
    // rom_array[16587] = 32'hFFFFFFF1;
    // rom_array[16588] = 32'hFFFFFFF1;
    // rom_array[16589] = 32'hFFFFFFF0;
    // rom_array[16590] = 32'hFFFFFFF0;
    // rom_array[16591] = 32'hFFFFFFF0;
    // rom_array[16592] = 32'hFFFFFFF0;
    // rom_array[16593] = 32'hFFFFFFF1;
    // rom_array[16594] = 32'hFFFFFFF1;
    // rom_array[16595] = 32'hFFFFFFF1;
    // rom_array[16596] = 32'hFFFFFFF1;
    // rom_array[16597] = 32'hFFFFFFF0;
    // rom_array[16598] = 32'hFFFFFFF0;
    // rom_array[16599] = 32'hFFFFFFF0;
    // rom_array[16600] = 32'hFFFFFFF0;
    // rom_array[16601] = 32'hFFFFFFF1;
    // rom_array[16602] = 32'hFFFFFFF1;
    // rom_array[16603] = 32'hFFFFFFF1;
    // rom_array[16604] = 32'hFFFFFFF1;
    // rom_array[16605] = 32'hFFFFFFF0;
    // rom_array[16606] = 32'hFFFFFFF0;
    // rom_array[16607] = 32'hFFFFFFF1;
    // rom_array[16608] = 32'hFFFFFFF1;
    // rom_array[16609] = 32'hFFFFFFF1;
    // rom_array[16610] = 32'hFFFFFFF1;
    // rom_array[16611] = 32'hFFFFFFF1;
    // rom_array[16612] = 32'hFFFFFFF1;
    // rom_array[16613] = 32'hFFFFFFF0;
    // rom_array[16614] = 32'hFFFFFFF0;
    // rom_array[16615] = 32'hFFFFFFF1;
    // rom_array[16616] = 32'hFFFFFFF1;
    // rom_array[16617] = 32'hFFFFFFF0;
    // rom_array[16618] = 32'hFFFFFFF0;
    // rom_array[16619] = 32'hFFFFFFF1;
    // rom_array[16620] = 32'hFFFFFFF1;
    // rom_array[16621] = 32'hFFFFFFF0;
    // rom_array[16622] = 32'hFFFFFFF0;
    // rom_array[16623] = 32'hFFFFFFF1;
    // rom_array[16624] = 32'hFFFFFFF1;
    // rom_array[16625] = 32'hFFFFFFF0;
    // rom_array[16626] = 32'hFFFFFFF0;
    // rom_array[16627] = 32'hFFFFFFF1;
    // rom_array[16628] = 32'hFFFFFFF1;
    // rom_array[16629] = 32'hFFFFFFF0;
    // rom_array[16630] = 32'hFFFFFFF0;
    // rom_array[16631] = 32'hFFFFFFF1;
    // rom_array[16632] = 32'hFFFFFFF1;
    // rom_array[16633] = 32'hFFFFFFF1;
    // rom_array[16634] = 32'hFFFFFFF1;
    // rom_array[16635] = 32'hFFFFFFF1;
    // rom_array[16636] = 32'hFFFFFFF1;
    // rom_array[16637] = 32'hFFFFFFF1;
    // rom_array[16638] = 32'hFFFFFFF1;
    // rom_array[16639] = 32'hFFFFFFF1;
    // rom_array[16640] = 32'hFFFFFFF1;
    // rom_array[16641] = 32'hFFFFFFF1;
    // rom_array[16642] = 32'hFFFFFFF1;
    // rom_array[16643] = 32'hFFFFFFF1;
    // rom_array[16644] = 32'hFFFFFFF1;
    // rom_array[16645] = 32'hFFFFFFF1;
    // rom_array[16646] = 32'hFFFFFFF1;
    // rom_array[16647] = 32'hFFFFFFF1;
    // rom_array[16648] = 32'hFFFFFFF1;
    // rom_array[16649] = 32'hFFFFFFF1;
    // rom_array[16650] = 32'hFFFFFFF1;
    // rom_array[16651] = 32'hFFFFFFF1;
    // rom_array[16652] = 32'hFFFFFFF1;
    // rom_array[16653] = 32'hFFFFFFF1;
    // rom_array[16654] = 32'hFFFFFFF1;
    // rom_array[16655] = 32'hFFFFFFF1;
    // rom_array[16656] = 32'hFFFFFFF1;
    // rom_array[16657] = 32'hFFFFFFF1;
    // rom_array[16658] = 32'hFFFFFFF1;
    // rom_array[16659] = 32'hFFFFFFF1;
    // rom_array[16660] = 32'hFFFFFFF1;
    // rom_array[16661] = 32'hFFFFFFF1;
    // rom_array[16662] = 32'hFFFFFFF1;
    // rom_array[16663] = 32'hFFFFFFF1;
    // rom_array[16664] = 32'hFFFFFFF1;
    // rom_array[16665] = 32'hFFFFFFF0;
    // rom_array[16666] = 32'hFFFFFFF0;
    // rom_array[16667] = 32'hFFFFFFF1;
    // rom_array[16668] = 32'hFFFFFFF1;
    // rom_array[16669] = 32'hFFFFFFF0;
    // rom_array[16670] = 32'hFFFFFFF0;
    // rom_array[16671] = 32'hFFFFFFF1;
    // rom_array[16672] = 32'hFFFFFFF1;
    // rom_array[16673] = 32'hFFFFFFF0;
    // rom_array[16674] = 32'hFFFFFFF0;
    // rom_array[16675] = 32'hFFFFFFF1;
    // rom_array[16676] = 32'hFFFFFFF1;
    // rom_array[16677] = 32'hFFFFFFF0;
    // rom_array[16678] = 32'hFFFFFFF0;
    // rom_array[16679] = 32'hFFFFFFF1;
    // rom_array[16680] = 32'hFFFFFFF1;
    // rom_array[16681] = 32'hFFFFFFF0;
    // rom_array[16682] = 32'hFFFFFFF0;
    // rom_array[16683] = 32'hFFFFFFF1;
    // rom_array[16684] = 32'hFFFFFFF1;
    // rom_array[16685] = 32'hFFFFFFF0;
    // rom_array[16686] = 32'hFFFFFFF0;
    // rom_array[16687] = 32'hFFFFFFF1;
    // rom_array[16688] = 32'hFFFFFFF1;
    // rom_array[16689] = 32'hFFFFFFF0;
    // rom_array[16690] = 32'hFFFFFFF0;
    // rom_array[16691] = 32'hFFFFFFF1;
    // rom_array[16692] = 32'hFFFFFFF1;
    // rom_array[16693] = 32'hFFFFFFF0;
    // rom_array[16694] = 32'hFFFFFFF0;
    // rom_array[16695] = 32'hFFFFFFF1;
    // rom_array[16696] = 32'hFFFFFFF1;
    // rom_array[16697] = 32'hFFFFFFF0;
    // rom_array[16698] = 32'hFFFFFFF0;
    // rom_array[16699] = 32'hFFFFFFF1;
    // rom_array[16700] = 32'hFFFFFFF1;
    // rom_array[16701] = 32'hFFFFFFF0;
    // rom_array[16702] = 32'hFFFFFFF0;
    // rom_array[16703] = 32'hFFFFFFF1;
    // rom_array[16704] = 32'hFFFFFFF1;
    // rom_array[16705] = 32'hFFFFFFF0;
    // rom_array[16706] = 32'hFFFFFFF0;
    // rom_array[16707] = 32'hFFFFFFF1;
    // rom_array[16708] = 32'hFFFFFFF1;
    // rom_array[16709] = 32'hFFFFFFF0;
    // rom_array[16710] = 32'hFFFFFFF0;
    // rom_array[16711] = 32'hFFFFFFF1;
    // rom_array[16712] = 32'hFFFFFFF1;
    // rom_array[16713] = 32'hFFFFFFF0;
    // rom_array[16714] = 32'hFFFFFFF0;
    // rom_array[16715] = 32'hFFFFFFF1;
    // rom_array[16716] = 32'hFFFFFFF1;
    // rom_array[16717] = 32'hFFFFFFF0;
    // rom_array[16718] = 32'hFFFFFFF0;
    // rom_array[16719] = 32'hFFFFFFF1;
    // rom_array[16720] = 32'hFFFFFFF1;
    // rom_array[16721] = 32'hFFFFFFF0;
    // rom_array[16722] = 32'hFFFFFFF0;
    // rom_array[16723] = 32'hFFFFFFF1;
    // rom_array[16724] = 32'hFFFFFFF1;
    // rom_array[16725] = 32'hFFFFFFF0;
    // rom_array[16726] = 32'hFFFFFFF0;
    // rom_array[16727] = 32'hFFFFFFF1;
    // rom_array[16728] = 32'hFFFFFFF1;
    // rom_array[16729] = 32'hFFFFFFF0;
    // rom_array[16730] = 32'hFFFFFFF0;
    // rom_array[16731] = 32'hFFFFFFF1;
    // rom_array[16732] = 32'hFFFFFFF1;
    // rom_array[16733] = 32'hFFFFFFF0;
    // rom_array[16734] = 32'hFFFFFFF0;
    // rom_array[16735] = 32'hFFFFFFF1;
    // rom_array[16736] = 32'hFFFFFFF1;
    // rom_array[16737] = 32'hFFFFFFF0;
    // rom_array[16738] = 32'hFFFFFFF0;
    // rom_array[16739] = 32'hFFFFFFF1;
    // rom_array[16740] = 32'hFFFFFFF1;
    // rom_array[16741] = 32'hFFFFFFF0;
    // rom_array[16742] = 32'hFFFFFFF0;
    // rom_array[16743] = 32'hFFFFFFF1;
    // rom_array[16744] = 32'hFFFFFFF1;
    // rom_array[16745] = 32'hFFFFFFF0;
    // rom_array[16746] = 32'hFFFFFFF0;
    // rom_array[16747] = 32'hFFFFFFF1;
    // rom_array[16748] = 32'hFFFFFFF1;
    // rom_array[16749] = 32'hFFFFFFF0;
    // rom_array[16750] = 32'hFFFFFFF0;
    // rom_array[16751] = 32'hFFFFFFF1;
    // rom_array[16752] = 32'hFFFFFFF1;
    // rom_array[16753] = 32'hFFFFFFF0;
    // rom_array[16754] = 32'hFFFFFFF0;
    // rom_array[16755] = 32'hFFFFFFF1;
    // rom_array[16756] = 32'hFFFFFFF1;
    // rom_array[16757] = 32'hFFFFFFF0;
    // rom_array[16758] = 32'hFFFFFFF0;
    // rom_array[16759] = 32'hFFFFFFF1;
    // rom_array[16760] = 32'hFFFFFFF1;
    // rom_array[16761] = 32'hFFFFFFF0;
    // rom_array[16762] = 32'hFFFFFFF0;
    // rom_array[16763] = 32'hFFFFFFF1;
    // rom_array[16764] = 32'hFFFFFFF1;
    // rom_array[16765] = 32'hFFFFFFF0;
    // rom_array[16766] = 32'hFFFFFFF0;
    // rom_array[16767] = 32'hFFFFFFF1;
    // rom_array[16768] = 32'hFFFFFFF1;
    // rom_array[16769] = 32'hFFFFFFF0;
    // rom_array[16770] = 32'hFFFFFFF0;
    // rom_array[16771] = 32'hFFFFFFF1;
    // rom_array[16772] = 32'hFFFFFFF1;
    // rom_array[16773] = 32'hFFFFFFF0;
    // rom_array[16774] = 32'hFFFFFFF0;
    // rom_array[16775] = 32'hFFFFFFF1;
    // rom_array[16776] = 32'hFFFFFFF1;
    // rom_array[16777] = 32'hFFFFFFF0;
    // rom_array[16778] = 32'hFFFFFFF0;
    // rom_array[16779] = 32'hFFFFFFF1;
    // rom_array[16780] = 32'hFFFFFFF1;
    // rom_array[16781] = 32'hFFFFFFF0;
    // rom_array[16782] = 32'hFFFFFFF0;
    // rom_array[16783] = 32'hFFFFFFF1;
    // rom_array[16784] = 32'hFFFFFFF1;
    // rom_array[16785] = 32'hFFFFFFF0;
    // rom_array[16786] = 32'hFFFFFFF0;
    // rom_array[16787] = 32'hFFFFFFF1;
    // rom_array[16788] = 32'hFFFFFFF1;
    // rom_array[16789] = 32'hFFFFFFF0;
    // rom_array[16790] = 32'hFFFFFFF0;
    // rom_array[16791] = 32'hFFFFFFF1;
    // rom_array[16792] = 32'hFFFFFFF1;
    // rom_array[16793] = 32'hFFFFFFF1;
    // rom_array[16794] = 32'hFFFFFFF1;
    // rom_array[16795] = 32'hFFFFFFF1;
    // rom_array[16796] = 32'hFFFFFFF1;
    // rom_array[16797] = 32'hFFFFFFF1;
    // rom_array[16798] = 32'hFFFFFFF1;
    // rom_array[16799] = 32'hFFFFFFF1;
    // rom_array[16800] = 32'hFFFFFFF1;
    // rom_array[16801] = 32'hFFFFFFF1;
    // rom_array[16802] = 32'hFFFFFFF1;
    // rom_array[16803] = 32'hFFFFFFF1;
    // rom_array[16804] = 32'hFFFFFFF1;
    // rom_array[16805] = 32'hFFFFFFF1;
    // rom_array[16806] = 32'hFFFFFFF1;
    // rom_array[16807] = 32'hFFFFFFF1;
    // rom_array[16808] = 32'hFFFFFFF1;
    // rom_array[16809] = 32'hFFFFFFF1;
    // rom_array[16810] = 32'hFFFFFFF1;
    // rom_array[16811] = 32'hFFFFFFF1;
    // rom_array[16812] = 32'hFFFFFFF1;
    // rom_array[16813] = 32'hFFFFFFF1;
    // rom_array[16814] = 32'hFFFFFFF1;
    // rom_array[16815] = 32'hFFFFFFF1;
    // rom_array[16816] = 32'hFFFFFFF1;
    // rom_array[16817] = 32'hFFFFFFF1;
    // rom_array[16818] = 32'hFFFFFFF1;
    // rom_array[16819] = 32'hFFFFFFF1;
    // rom_array[16820] = 32'hFFFFFFF1;
    // rom_array[16821] = 32'hFFFFFFF1;
    // rom_array[16822] = 32'hFFFFFFF1;
    // rom_array[16823] = 32'hFFFFFFF1;
    // rom_array[16824] = 32'hFFFFFFF1;
    // rom_array[16825] = 32'hFFFFFFF1;
    // rom_array[16826] = 32'hFFFFFFF1;
    // rom_array[16827] = 32'hFFFFFFF1;
    // rom_array[16828] = 32'hFFFFFFF1;
    // rom_array[16829] = 32'hFFFFFFF1;
    // rom_array[16830] = 32'hFFFFFFF1;
    // rom_array[16831] = 32'hFFFFFFF1;
    // rom_array[16832] = 32'hFFFFFFF1;
    // rom_array[16833] = 32'hFFFFFFF1;
    // rom_array[16834] = 32'hFFFFFFF1;
    // rom_array[16835] = 32'hFFFFFFF1;
    // rom_array[16836] = 32'hFFFFFFF1;
    // rom_array[16837] = 32'hFFFFFFF1;
    // rom_array[16838] = 32'hFFFFFFF1;
    // rom_array[16839] = 32'hFFFFFFF1;
    // rom_array[16840] = 32'hFFFFFFF1;
    // rom_array[16841] = 32'hFFFFFFF1;
    // rom_array[16842] = 32'hFFFFFFF1;
    // rom_array[16843] = 32'hFFFFFFF1;
    // rom_array[16844] = 32'hFFFFFFF1;
    // rom_array[16845] = 32'hFFFFFFF1;
    // rom_array[16846] = 32'hFFFFFFF1;
    // rom_array[16847] = 32'hFFFFFFF1;
    // rom_array[16848] = 32'hFFFFFFF1;
    // rom_array[16849] = 32'hFFFFFFF1;
    // rom_array[16850] = 32'hFFFFFFF1;
    // rom_array[16851] = 32'hFFFFFFF1;
    // rom_array[16852] = 32'hFFFFFFF1;
    // rom_array[16853] = 32'hFFFFFFF1;
    // rom_array[16854] = 32'hFFFFFFF1;
    // rom_array[16855] = 32'hFFFFFFF1;
    // rom_array[16856] = 32'hFFFFFFF1;
    // rom_array[16857] = 32'hFFFFFFF0;
    // rom_array[16858] = 32'hFFFFFFF0;
    // rom_array[16859] = 32'hFFFFFFF1;
    // rom_array[16860] = 32'hFFFFFFF1;
    // rom_array[16861] = 32'hFFFFFFF0;
    // rom_array[16862] = 32'hFFFFFFF0;
    // rom_array[16863] = 32'hFFFFFFF1;
    // rom_array[16864] = 32'hFFFFFFF1;
    // rom_array[16865] = 32'hFFFFFFF0;
    // rom_array[16866] = 32'hFFFFFFF0;
    // rom_array[16867] = 32'hFFFFFFF1;
    // rom_array[16868] = 32'hFFFFFFF1;
    // rom_array[16869] = 32'hFFFFFFF0;
    // rom_array[16870] = 32'hFFFFFFF0;
    // rom_array[16871] = 32'hFFFFFFF1;
    // rom_array[16872] = 32'hFFFFFFF1;
    // rom_array[16873] = 32'hFFFFFFF0;
    // rom_array[16874] = 32'hFFFFFFF0;
    // rom_array[16875] = 32'hFFFFFFF1;
    // rom_array[16876] = 32'hFFFFFFF1;
    // rom_array[16877] = 32'hFFFFFFF0;
    // rom_array[16878] = 32'hFFFFFFF0;
    // rom_array[16879] = 32'hFFFFFFF1;
    // rom_array[16880] = 32'hFFFFFFF1;
    // rom_array[16881] = 32'hFFFFFFF0;
    // rom_array[16882] = 32'hFFFFFFF0;
    // rom_array[16883] = 32'hFFFFFFF1;
    // rom_array[16884] = 32'hFFFFFFF1;
    // rom_array[16885] = 32'hFFFFFFF0;
    // rom_array[16886] = 32'hFFFFFFF0;
    // rom_array[16887] = 32'hFFFFFFF1;
    // rom_array[16888] = 32'hFFFFFFF1;
    // rom_array[16889] = 32'hFFFFFFF0;
    // rom_array[16890] = 32'hFFFFFFF0;
    // rom_array[16891] = 32'hFFFFFFF1;
    // rom_array[16892] = 32'hFFFFFFF1;
    // rom_array[16893] = 32'hFFFFFFF0;
    // rom_array[16894] = 32'hFFFFFFF0;
    // rom_array[16895] = 32'hFFFFFFF1;
    // rom_array[16896] = 32'hFFFFFFF1;
    // rom_array[16897] = 32'hFFFFFFF0;
    // rom_array[16898] = 32'hFFFFFFF0;
    // rom_array[16899] = 32'hFFFFFFF1;
    // rom_array[16900] = 32'hFFFFFFF1;
    // rom_array[16901] = 32'hFFFFFFF0;
    // rom_array[16902] = 32'hFFFFFFF0;
    // rom_array[16903] = 32'hFFFFFFF1;
    // rom_array[16904] = 32'hFFFFFFF1;
    // rom_array[16905] = 32'hFFFFFFF0;
    // rom_array[16906] = 32'hFFFFFFF0;
    // rom_array[16907] = 32'hFFFFFFF1;
    // rom_array[16908] = 32'hFFFFFFF1;
    // rom_array[16909] = 32'hFFFFFFF0;
    // rom_array[16910] = 32'hFFFFFFF0;
    // rom_array[16911] = 32'hFFFFFFF1;
    // rom_array[16912] = 32'hFFFFFFF1;
    // rom_array[16913] = 32'hFFFFFFF0;
    // rom_array[16914] = 32'hFFFFFFF0;
    // rom_array[16915] = 32'hFFFFFFF1;
    // rom_array[16916] = 32'hFFFFFFF1;
    // rom_array[16917] = 32'hFFFFFFF0;
    // rom_array[16918] = 32'hFFFFFFF0;
    // rom_array[16919] = 32'hFFFFFFF1;
    // rom_array[16920] = 32'hFFFFFFF1;
    // rom_array[16921] = 32'hFFFFFFF1;
    // rom_array[16922] = 32'hFFFFFFF1;
    // rom_array[16923] = 32'hFFFFFFF1;
    // rom_array[16924] = 32'hFFFFFFF1;
    // rom_array[16925] = 32'hFFFFFFF1;
    // rom_array[16926] = 32'hFFFFFFF1;
    // rom_array[16927] = 32'hFFFFFFF1;
    // rom_array[16928] = 32'hFFFFFFF1;
    // rom_array[16929] = 32'hFFFFFFF1;
    // rom_array[16930] = 32'hFFFFFFF1;
    // rom_array[16931] = 32'hFFFFFFF1;
    // rom_array[16932] = 32'hFFFFFFF1;
    // rom_array[16933] = 32'hFFFFFFF1;
    // rom_array[16934] = 32'hFFFFFFF1;
    // rom_array[16935] = 32'hFFFFFFF1;
    // rom_array[16936] = 32'hFFFFFFF1;
    // rom_array[16937] = 32'hFFFFFFF1;
    // rom_array[16938] = 32'hFFFFFFF1;
    // rom_array[16939] = 32'hFFFFFFF1;
    // rom_array[16940] = 32'hFFFFFFF1;
    // rom_array[16941] = 32'hFFFFFFF1;
    // rom_array[16942] = 32'hFFFFFFF1;
    // rom_array[16943] = 32'hFFFFFFF1;
    // rom_array[16944] = 32'hFFFFFFF1;
    // rom_array[16945] = 32'hFFFFFFF1;
    // rom_array[16946] = 32'hFFFFFFF1;
    // rom_array[16947] = 32'hFFFFFFF1;
    // rom_array[16948] = 32'hFFFFFFF1;
    // rom_array[16949] = 32'hFFFFFFF1;
    // rom_array[16950] = 32'hFFFFFFF1;
    // rom_array[16951] = 32'hFFFFFFF1;
    // rom_array[16952] = 32'hFFFFFFF1;
    // rom_array[16953] = 32'hFFFFFFF1;
    // rom_array[16954] = 32'hFFFFFFF1;
    // rom_array[16955] = 32'hFFFFFFF1;
    // rom_array[16956] = 32'hFFFFFFF1;
    // rom_array[16957] = 32'hFFFFFFF1;
    // rom_array[16958] = 32'hFFFFFFF1;
    // rom_array[16959] = 32'hFFFFFFF1;
    // rom_array[16960] = 32'hFFFFFFF1;
    // rom_array[16961] = 32'hFFFFFFF1;
    // rom_array[16962] = 32'hFFFFFFF1;
    // rom_array[16963] = 32'hFFFFFFF1;
    // rom_array[16964] = 32'hFFFFFFF1;
    // rom_array[16965] = 32'hFFFFFFF1;
    // rom_array[16966] = 32'hFFFFFFF1;
    // rom_array[16967] = 32'hFFFFFFF1;
    // rom_array[16968] = 32'hFFFFFFF1;
    // rom_array[16969] = 32'hFFFFFFF1;
    // rom_array[16970] = 32'hFFFFFFF1;
    // rom_array[16971] = 32'hFFFFFFF1;
    // rom_array[16972] = 32'hFFFFFFF1;
    // rom_array[16973] = 32'hFFFFFFF1;
    // rom_array[16974] = 32'hFFFFFFF1;
    // rom_array[16975] = 32'hFFFFFFF1;
    // rom_array[16976] = 32'hFFFFFFF1;
    // rom_array[16977] = 32'hFFFFFFF1;
    // rom_array[16978] = 32'hFFFFFFF1;
    // rom_array[16979] = 32'hFFFFFFF1;
    // rom_array[16980] = 32'hFFFFFFF1;
    // rom_array[16981] = 32'hFFFFFFF1;
    // rom_array[16982] = 32'hFFFFFFF1;
    // rom_array[16983] = 32'hFFFFFFF1;
    // rom_array[16984] = 32'hFFFFFFF1;
    // rom_array[16985] = 32'hFFFFFFF0;
    // rom_array[16986] = 32'hFFFFFFF0;
    // rom_array[16987] = 32'hFFFFFFF1;
    // rom_array[16988] = 32'hFFFFFFF1;
    // rom_array[16989] = 32'hFFFFFFF0;
    // rom_array[16990] = 32'hFFFFFFF0;
    // rom_array[16991] = 32'hFFFFFFF1;
    // rom_array[16992] = 32'hFFFFFFF1;
    // rom_array[16993] = 32'hFFFFFFF0;
    // rom_array[16994] = 32'hFFFFFFF0;
    // rom_array[16995] = 32'hFFFFFFF1;
    // rom_array[16996] = 32'hFFFFFFF1;
    // rom_array[16997] = 32'hFFFFFFF0;
    // rom_array[16998] = 32'hFFFFFFF0;
    // rom_array[16999] = 32'hFFFFFFF1;
    // rom_array[17000] = 32'hFFFFFFF1;
    // rom_array[17001] = 32'hFFFFFFF0;
    // rom_array[17002] = 32'hFFFFFFF0;
    // rom_array[17003] = 32'hFFFFFFF1;
    // rom_array[17004] = 32'hFFFFFFF1;
    // rom_array[17005] = 32'hFFFFFFF0;
    // rom_array[17006] = 32'hFFFFFFF0;
    // rom_array[17007] = 32'hFFFFFFF1;
    // rom_array[17008] = 32'hFFFFFFF1;
    // rom_array[17009] = 32'hFFFFFFF0;
    // rom_array[17010] = 32'hFFFFFFF0;
    // rom_array[17011] = 32'hFFFFFFF1;
    // rom_array[17012] = 32'hFFFFFFF1;
    // rom_array[17013] = 32'hFFFFFFF0;
    // rom_array[17014] = 32'hFFFFFFF0;
    // rom_array[17015] = 32'hFFFFFFF1;
    // rom_array[17016] = 32'hFFFFFFF1;
    // rom_array[17017] = 32'hFFFFFFF0;
    // rom_array[17018] = 32'hFFFFFFF0;
    // rom_array[17019] = 32'hFFFFFFF1;
    // rom_array[17020] = 32'hFFFFFFF1;
    // rom_array[17021] = 32'hFFFFFFF0;
    // rom_array[17022] = 32'hFFFFFFF0;
    // rom_array[17023] = 32'hFFFFFFF1;
    // rom_array[17024] = 32'hFFFFFFF1;
    // rom_array[17025] = 32'hFFFFFFF0;
    // rom_array[17026] = 32'hFFFFFFF0;
    // rom_array[17027] = 32'hFFFFFFF1;
    // rom_array[17028] = 32'hFFFFFFF1;
    // rom_array[17029] = 32'hFFFFFFF0;
    // rom_array[17030] = 32'hFFFFFFF0;
    // rom_array[17031] = 32'hFFFFFFF1;
    // rom_array[17032] = 32'hFFFFFFF1;
    // rom_array[17033] = 32'hFFFFFFF0;
    // rom_array[17034] = 32'hFFFFFFF0;
    // rom_array[17035] = 32'hFFFFFFF1;
    // rom_array[17036] = 32'hFFFFFFF1;
    // rom_array[17037] = 32'hFFFFFFF0;
    // rom_array[17038] = 32'hFFFFFFF0;
    // rom_array[17039] = 32'hFFFFFFF1;
    // rom_array[17040] = 32'hFFFFFFF1;
    // rom_array[17041] = 32'hFFFFFFF0;
    // rom_array[17042] = 32'hFFFFFFF0;
    // rom_array[17043] = 32'hFFFFFFF1;
    // rom_array[17044] = 32'hFFFFFFF1;
    // rom_array[17045] = 32'hFFFFFFF0;
    // rom_array[17046] = 32'hFFFFFFF0;
    // rom_array[17047] = 32'hFFFFFFF1;
    // rom_array[17048] = 32'hFFFFFFF1;
    // rom_array[17049] = 32'hFFFFFFF0;
    // rom_array[17050] = 32'hFFFFFFF0;
    // rom_array[17051] = 32'hFFFFFFF0;
    // rom_array[17052] = 32'hFFFFFFF0;
    // rom_array[17053] = 32'hFFFFFFF0;
    // rom_array[17054] = 32'hFFFFFFF0;
    // rom_array[17055] = 32'hFFFFFFF1;
    // rom_array[17056] = 32'hFFFFFFF1;
    // rom_array[17057] = 32'hFFFFFFF0;
    // rom_array[17058] = 32'hFFFFFFF0;
    // rom_array[17059] = 32'hFFFFFFF0;
    // rom_array[17060] = 32'hFFFFFFF0;
    // rom_array[17061] = 32'hFFFFFFF0;
    // rom_array[17062] = 32'hFFFFFFF0;
    // rom_array[17063] = 32'hFFFFFFF1;
    // rom_array[17064] = 32'hFFFFFFF1;
    // rom_array[17065] = 32'hFFFFFFF0;
    // rom_array[17066] = 32'hFFFFFFF0;
    // rom_array[17067] = 32'hFFFFFFF0;
    // rom_array[17068] = 32'hFFFFFFF0;
    // rom_array[17069] = 32'hFFFFFFF1;
    // rom_array[17070] = 32'hFFFFFFF1;
    // rom_array[17071] = 32'hFFFFFFF1;
    // rom_array[17072] = 32'hFFFFFFF1;
    // rom_array[17073] = 32'hFFFFFFF0;
    // rom_array[17074] = 32'hFFFFFFF0;
    // rom_array[17075] = 32'hFFFFFFF0;
    // rom_array[17076] = 32'hFFFFFFF0;
    // rom_array[17077] = 32'hFFFFFFF1;
    // rom_array[17078] = 32'hFFFFFFF1;
    // rom_array[17079] = 32'hFFFFFFF1;
    // rom_array[17080] = 32'hFFFFFFF1;
    // rom_array[17081] = 32'hFFFFFFF0;
    // rom_array[17082] = 32'hFFFFFFF0;
    // rom_array[17083] = 32'hFFFFFFF0;
    // rom_array[17084] = 32'hFFFFFFF0;
    // rom_array[17085] = 32'hFFFFFFF1;
    // rom_array[17086] = 32'hFFFFFFF1;
    // rom_array[17087] = 32'hFFFFFFF1;
    // rom_array[17088] = 32'hFFFFFFF1;
    // rom_array[17089] = 32'hFFFFFFF0;
    // rom_array[17090] = 32'hFFFFFFF0;
    // rom_array[17091] = 32'hFFFFFFF0;
    // rom_array[17092] = 32'hFFFFFFF0;
    // rom_array[17093] = 32'hFFFFFFF1;
    // rom_array[17094] = 32'hFFFFFFF1;
    // rom_array[17095] = 32'hFFFFFFF1;
    // rom_array[17096] = 32'hFFFFFFF1;
    // rom_array[17097] = 32'hFFFFFFF0;
    // rom_array[17098] = 32'hFFFFFFF0;
    // rom_array[17099] = 32'hFFFFFFF0;
    // rom_array[17100] = 32'hFFFFFFF0;
    // rom_array[17101] = 32'hFFFFFFF1;
    // rom_array[17102] = 32'hFFFFFFF1;
    // rom_array[17103] = 32'hFFFFFFF1;
    // rom_array[17104] = 32'hFFFFFFF1;
    // rom_array[17105] = 32'hFFFFFFF0;
    // rom_array[17106] = 32'hFFFFFFF0;
    // rom_array[17107] = 32'hFFFFFFF0;
    // rom_array[17108] = 32'hFFFFFFF0;
    // rom_array[17109] = 32'hFFFFFFF1;
    // rom_array[17110] = 32'hFFFFFFF1;
    // rom_array[17111] = 32'hFFFFFFF1;
    // rom_array[17112] = 32'hFFFFFFF1;
    // rom_array[17113] = 32'hFFFFFFF0;
    // rom_array[17114] = 32'hFFFFFFF0;
    // rom_array[17115] = 32'hFFFFFFF1;
    // rom_array[17116] = 32'hFFFFFFF1;
    // rom_array[17117] = 32'hFFFFFFF0;
    // rom_array[17118] = 32'hFFFFFFF0;
    // rom_array[17119] = 32'hFFFFFFF1;
    // rom_array[17120] = 32'hFFFFFFF1;
    // rom_array[17121] = 32'hFFFFFFF0;
    // rom_array[17122] = 32'hFFFFFFF0;
    // rom_array[17123] = 32'hFFFFFFF1;
    // rom_array[17124] = 32'hFFFFFFF1;
    // rom_array[17125] = 32'hFFFFFFF0;
    // rom_array[17126] = 32'hFFFFFFF0;
    // rom_array[17127] = 32'hFFFFFFF1;
    // rom_array[17128] = 32'hFFFFFFF1;
    // rom_array[17129] = 32'hFFFFFFF0;
    // rom_array[17130] = 32'hFFFFFFF0;
    // rom_array[17131] = 32'hFFFFFFF1;
    // rom_array[17132] = 32'hFFFFFFF1;
    // rom_array[17133] = 32'hFFFFFFF0;
    // rom_array[17134] = 32'hFFFFFFF0;
    // rom_array[17135] = 32'hFFFFFFF1;
    // rom_array[17136] = 32'hFFFFFFF1;
    // rom_array[17137] = 32'hFFFFFFF0;
    // rom_array[17138] = 32'hFFFFFFF0;
    // rom_array[17139] = 32'hFFFFFFF1;
    // rom_array[17140] = 32'hFFFFFFF1;
    // rom_array[17141] = 32'hFFFFFFF0;
    // rom_array[17142] = 32'hFFFFFFF0;
    // rom_array[17143] = 32'hFFFFFFF1;
    // rom_array[17144] = 32'hFFFFFFF1;
    // rom_array[17145] = 32'hFFFFFFF0;
    // rom_array[17146] = 32'hFFFFFFF0;
    // rom_array[17147] = 32'hFFFFFFF0;
    // rom_array[17148] = 32'hFFFFFFF0;
    // rom_array[17149] = 32'hFFFFFFF1;
    // rom_array[17150] = 32'hFFFFFFF1;
    // rom_array[17151] = 32'hFFFFFFF1;
    // rom_array[17152] = 32'hFFFFFFF1;
    // rom_array[17153] = 32'hFFFFFFF0;
    // rom_array[17154] = 32'hFFFFFFF0;
    // rom_array[17155] = 32'hFFFFFFF0;
    // rom_array[17156] = 32'hFFFFFFF0;
    // rom_array[17157] = 32'hFFFFFFF1;
    // rom_array[17158] = 32'hFFFFFFF1;
    // rom_array[17159] = 32'hFFFFFFF1;
    // rom_array[17160] = 32'hFFFFFFF1;
    // rom_array[17161] = 32'hFFFFFFF1;
    // rom_array[17162] = 32'hFFFFFFF1;
    // rom_array[17163] = 32'hFFFFFFF1;
    // rom_array[17164] = 32'hFFFFFFF1;
    // rom_array[17165] = 32'hFFFFFFF1;
    // rom_array[17166] = 32'hFFFFFFF1;
    // rom_array[17167] = 32'hFFFFFFF1;
    // rom_array[17168] = 32'hFFFFFFF1;
    // rom_array[17169] = 32'hFFFFFFF1;
    // rom_array[17170] = 32'hFFFFFFF1;
    // rom_array[17171] = 32'hFFFFFFF1;
    // rom_array[17172] = 32'hFFFFFFF1;
    // rom_array[17173] = 32'hFFFFFFF1;
    // rom_array[17174] = 32'hFFFFFFF1;
    // rom_array[17175] = 32'hFFFFFFF1;
    // rom_array[17176] = 32'hFFFFFFF1;
    // rom_array[17177] = 32'hFFFFFFF1;
    // rom_array[17178] = 32'hFFFFFFF1;
    // rom_array[17179] = 32'hFFFFFFF1;
    // rom_array[17180] = 32'hFFFFFFF1;
    // rom_array[17181] = 32'hFFFFFFF1;
    // rom_array[17182] = 32'hFFFFFFF1;
    // rom_array[17183] = 32'hFFFFFFF1;
    // rom_array[17184] = 32'hFFFFFFF1;
    // rom_array[17185] = 32'hFFFFFFF1;
    // rom_array[17186] = 32'hFFFFFFF1;
    // rom_array[17187] = 32'hFFFFFFF1;
    // rom_array[17188] = 32'hFFFFFFF1;
    // rom_array[17189] = 32'hFFFFFFF1;
    // rom_array[17190] = 32'hFFFFFFF1;
    // rom_array[17191] = 32'hFFFFFFF1;
    // rom_array[17192] = 32'hFFFFFFF1;
    // rom_array[17193] = 32'hFFFFFFF0;
    // rom_array[17194] = 32'hFFFFFFF0;
    // rom_array[17195] = 32'hFFFFFFF1;
    // rom_array[17196] = 32'hFFFFFFF1;
    // rom_array[17197] = 32'hFFFFFFF0;
    // rom_array[17198] = 32'hFFFFFFF0;
    // rom_array[17199] = 32'hFFFFFFF1;
    // rom_array[17200] = 32'hFFFFFFF1;
    // rom_array[17201] = 32'hFFFFFFF0;
    // rom_array[17202] = 32'hFFFFFFF0;
    // rom_array[17203] = 32'hFFFFFFF1;
    // rom_array[17204] = 32'hFFFFFFF1;
    // rom_array[17205] = 32'hFFFFFFF0;
    // rom_array[17206] = 32'hFFFFFFF0;
    // rom_array[17207] = 32'hFFFFFFF1;
    // rom_array[17208] = 32'hFFFFFFF1;
    // rom_array[17209] = 32'hFFFFFFF0;
    // rom_array[17210] = 32'hFFFFFFF0;
    // rom_array[17211] = 32'hFFFFFFF1;
    // rom_array[17212] = 32'hFFFFFFF1;
    // rom_array[17213] = 32'hFFFFFFF0;
    // rom_array[17214] = 32'hFFFFFFF0;
    // rom_array[17215] = 32'hFFFFFFF1;
    // rom_array[17216] = 32'hFFFFFFF1;
    // rom_array[17217] = 32'hFFFFFFF0;
    // rom_array[17218] = 32'hFFFFFFF0;
    // rom_array[17219] = 32'hFFFFFFF1;
    // rom_array[17220] = 32'hFFFFFFF1;
    // rom_array[17221] = 32'hFFFFFFF0;
    // rom_array[17222] = 32'hFFFFFFF0;
    // rom_array[17223] = 32'hFFFFFFF1;
    // rom_array[17224] = 32'hFFFFFFF1;
    // rom_array[17225] = 32'hFFFFFFF0;
    // rom_array[17226] = 32'hFFFFFFF0;
    // rom_array[17227] = 32'hFFFFFFF1;
    // rom_array[17228] = 32'hFFFFFFF1;
    // rom_array[17229] = 32'hFFFFFFF0;
    // rom_array[17230] = 32'hFFFFFFF0;
    // rom_array[17231] = 32'hFFFFFFF1;
    // rom_array[17232] = 32'hFFFFFFF1;
    // rom_array[17233] = 32'hFFFFFFF0;
    // rom_array[17234] = 32'hFFFFFFF0;
    // rom_array[17235] = 32'hFFFFFFF1;
    // rom_array[17236] = 32'hFFFFFFF1;
    // rom_array[17237] = 32'hFFFFFFF0;
    // rom_array[17238] = 32'hFFFFFFF0;
    // rom_array[17239] = 32'hFFFFFFF1;
    // rom_array[17240] = 32'hFFFFFFF1;
    // rom_array[17241] = 32'hFFFFFFF0;
    // rom_array[17242] = 32'hFFFFFFF0;
    // rom_array[17243] = 32'hFFFFFFF1;
    // rom_array[17244] = 32'hFFFFFFF1;
    // rom_array[17245] = 32'hFFFFFFF0;
    // rom_array[17246] = 32'hFFFFFFF0;
    // rom_array[17247] = 32'hFFFFFFF1;
    // rom_array[17248] = 32'hFFFFFFF1;
    // rom_array[17249] = 32'hFFFFFFF0;
    // rom_array[17250] = 32'hFFFFFFF0;
    // rom_array[17251] = 32'hFFFFFFF1;
    // rom_array[17252] = 32'hFFFFFFF1;
    // rom_array[17253] = 32'hFFFFFFF0;
    // rom_array[17254] = 32'hFFFFFFF0;
    // rom_array[17255] = 32'hFFFFFFF1;
    // rom_array[17256] = 32'hFFFFFFF1;
    // rom_array[17257] = 32'hFFFFFFF0;
    // rom_array[17258] = 32'hFFFFFFF0;
    // rom_array[17259] = 32'hFFFFFFF1;
    // rom_array[17260] = 32'hFFFFFFF1;
    // rom_array[17261] = 32'hFFFFFFF0;
    // rom_array[17262] = 32'hFFFFFFF0;
    // rom_array[17263] = 32'hFFFFFFF1;
    // rom_array[17264] = 32'hFFFFFFF1;
    // rom_array[17265] = 32'hFFFFFFF0;
    // rom_array[17266] = 32'hFFFFFFF0;
    // rom_array[17267] = 32'hFFFFFFF1;
    // rom_array[17268] = 32'hFFFFFFF1;
    // rom_array[17269] = 32'hFFFFFFF0;
    // rom_array[17270] = 32'hFFFFFFF0;
    // rom_array[17271] = 32'hFFFFFFF1;
    // rom_array[17272] = 32'hFFFFFFF1;
    // rom_array[17273] = 32'hFFFFFFF0;
    // rom_array[17274] = 32'hFFFFFFF0;
    // rom_array[17275] = 32'hFFFFFFF1;
    // rom_array[17276] = 32'hFFFFFFF1;
    // rom_array[17277] = 32'hFFFFFFF0;
    // rom_array[17278] = 32'hFFFFFFF0;
    // rom_array[17279] = 32'hFFFFFFF1;
    // rom_array[17280] = 32'hFFFFFFF1;
    // rom_array[17281] = 32'hFFFFFFF0;
    // rom_array[17282] = 32'hFFFFFFF0;
    // rom_array[17283] = 32'hFFFFFFF1;
    // rom_array[17284] = 32'hFFFFFFF1;
    // rom_array[17285] = 32'hFFFFFFF0;
    // rom_array[17286] = 32'hFFFFFFF0;
    // rom_array[17287] = 32'hFFFFFFF1;
    // rom_array[17288] = 32'hFFFFFFF1;
    // rom_array[17289] = 32'hFFFFFFF0;
    // rom_array[17290] = 32'hFFFFFFF0;
    // rom_array[17291] = 32'hFFFFFFF1;
    // rom_array[17292] = 32'hFFFFFFF1;
    // rom_array[17293] = 32'hFFFFFFF0;
    // rom_array[17294] = 32'hFFFFFFF0;
    // rom_array[17295] = 32'hFFFFFFF1;
    // rom_array[17296] = 32'hFFFFFFF1;
    // rom_array[17297] = 32'hFFFFFFF0;
    // rom_array[17298] = 32'hFFFFFFF0;
    // rom_array[17299] = 32'hFFFFFFF1;
    // rom_array[17300] = 32'hFFFFFFF1;
    // rom_array[17301] = 32'hFFFFFFF0;
    // rom_array[17302] = 32'hFFFFFFF0;
    // rom_array[17303] = 32'hFFFFFFF1;
    // rom_array[17304] = 32'hFFFFFFF1;
    // rom_array[17305] = 32'hFFFFFFF0;
    // rom_array[17306] = 32'hFFFFFFF0;
    // rom_array[17307] = 32'hFFFFFFF1;
    // rom_array[17308] = 32'hFFFFFFF1;
    // rom_array[17309] = 32'hFFFFFFF0;
    // rom_array[17310] = 32'hFFFFFFF0;
    // rom_array[17311] = 32'hFFFFFFF1;
    // rom_array[17312] = 32'hFFFFFFF1;
    // rom_array[17313] = 32'hFFFFFFF0;
    // rom_array[17314] = 32'hFFFFFFF0;
    // rom_array[17315] = 32'hFFFFFFF1;
    // rom_array[17316] = 32'hFFFFFFF1;
    // rom_array[17317] = 32'hFFFFFFF0;
    // rom_array[17318] = 32'hFFFFFFF0;
    // rom_array[17319] = 32'hFFFFFFF1;
    // rom_array[17320] = 32'hFFFFFFF1;
    // rom_array[17321] = 32'hFFFFFFF1;
    // rom_array[17322] = 32'hFFFFFFF1;
    // rom_array[17323] = 32'hFFFFFFF1;
    // rom_array[17324] = 32'hFFFFFFF1;
    // rom_array[17325] = 32'hFFFFFFF1;
    // rom_array[17326] = 32'hFFFFFFF1;
    // rom_array[17327] = 32'hFFFFFFF1;
    // rom_array[17328] = 32'hFFFFFFF1;
    // rom_array[17329] = 32'hFFFFFFF1;
    // rom_array[17330] = 32'hFFFFFFF1;
    // rom_array[17331] = 32'hFFFFFFF1;
    // rom_array[17332] = 32'hFFFFFFF1;
    // rom_array[17333] = 32'hFFFFFFF1;
    // rom_array[17334] = 32'hFFFFFFF1;
    // rom_array[17335] = 32'hFFFFFFF1;
    // rom_array[17336] = 32'hFFFFFFF1;
    // rom_array[17337] = 32'hFFFFFFF1;
    // rom_array[17338] = 32'hFFFFFFF1;
    // rom_array[17339] = 32'hFFFFFFF1;
    // rom_array[17340] = 32'hFFFFFFF1;
    // rom_array[17341] = 32'hFFFFFFF1;
    // rom_array[17342] = 32'hFFFFFFF1;
    // rom_array[17343] = 32'hFFFFFFF1;
    // rom_array[17344] = 32'hFFFFFFF1;
    // rom_array[17345] = 32'hFFFFFFF1;
    // rom_array[17346] = 32'hFFFFFFF1;
    // rom_array[17347] = 32'hFFFFFFF1;
    // rom_array[17348] = 32'hFFFFFFF1;
    // rom_array[17349] = 32'hFFFFFFF1;
    // rom_array[17350] = 32'hFFFFFFF1;
    // rom_array[17351] = 32'hFFFFFFF1;
    // rom_array[17352] = 32'hFFFFFFF1;
    // rom_array[17353] = 32'hFFFFFFF1;
    // rom_array[17354] = 32'hFFFFFFF1;
    // rom_array[17355] = 32'hFFFFFFF1;
    // rom_array[17356] = 32'hFFFFFFF1;
    // rom_array[17357] = 32'hFFFFFFF1;
    // rom_array[17358] = 32'hFFFFFFF1;
    // rom_array[17359] = 32'hFFFFFFF1;
    // rom_array[17360] = 32'hFFFFFFF1;
    // rom_array[17361] = 32'hFFFFFFF1;
    // rom_array[17362] = 32'hFFFFFFF1;
    // rom_array[17363] = 32'hFFFFFFF1;
    // rom_array[17364] = 32'hFFFFFFF1;
    // rom_array[17365] = 32'hFFFFFFF1;
    // rom_array[17366] = 32'hFFFFFFF1;
    // rom_array[17367] = 32'hFFFFFFF1;
    // rom_array[17368] = 32'hFFFFFFF1;
    // rom_array[17369] = 32'hFFFFFFF0;
    // rom_array[17370] = 32'hFFFFFFF0;
    // rom_array[17371] = 32'hFFFFFFF0;
    // rom_array[17372] = 32'hFFFFFFF0;
    // rom_array[17373] = 32'hFFFFFFF1;
    // rom_array[17374] = 32'hFFFFFFF1;
    // rom_array[17375] = 32'hFFFFFFF1;
    // rom_array[17376] = 32'hFFFFFFF1;
    // rom_array[17377] = 32'hFFFFFFF0;
    // rom_array[17378] = 32'hFFFFFFF0;
    // rom_array[17379] = 32'hFFFFFFF0;
    // rom_array[17380] = 32'hFFFFFFF0;
    // rom_array[17381] = 32'hFFFFFFF1;
    // rom_array[17382] = 32'hFFFFFFF1;
    // rom_array[17383] = 32'hFFFFFFF1;
    // rom_array[17384] = 32'hFFFFFFF1;
    // rom_array[17385] = 32'hFFFFFFF1;
    // rom_array[17386] = 32'hFFFFFFF1;
    // rom_array[17387] = 32'hFFFFFFF1;
    // rom_array[17388] = 32'hFFFFFFF1;
    // rom_array[17389] = 32'hFFFFFFF1;
    // rom_array[17390] = 32'hFFFFFFF1;
    // rom_array[17391] = 32'hFFFFFFF1;
    // rom_array[17392] = 32'hFFFFFFF1;
    // rom_array[17393] = 32'hFFFFFFF1;
    // rom_array[17394] = 32'hFFFFFFF1;
    // rom_array[17395] = 32'hFFFFFFF1;
    // rom_array[17396] = 32'hFFFFFFF1;
    // rom_array[17397] = 32'hFFFFFFF1;
    // rom_array[17398] = 32'hFFFFFFF1;
    // rom_array[17399] = 32'hFFFFFFF1;
    // rom_array[17400] = 32'hFFFFFFF1;
    // rom_array[17401] = 32'hFFFFFFF0;
    // rom_array[17402] = 32'hFFFFFFF0;
    // rom_array[17403] = 32'hFFFFFFF0;
    // rom_array[17404] = 32'hFFFFFFF0;
    // rom_array[17405] = 32'hFFFFFFF1;
    // rom_array[17406] = 32'hFFFFFFF1;
    // rom_array[17407] = 32'hFFFFFFF1;
    // rom_array[17408] = 32'hFFFFFFF1;
    // rom_array[17409] = 32'hFFFFFFF0;
    // rom_array[17410] = 32'hFFFFFFF0;
    // rom_array[17411] = 32'hFFFFFFF0;
    // rom_array[17412] = 32'hFFFFFFF0;
    // rom_array[17413] = 32'hFFFFFFF1;
    // rom_array[17414] = 32'hFFFFFFF1;
    // rom_array[17415] = 32'hFFFFFFF1;
    // rom_array[17416] = 32'hFFFFFFF1;
    // rom_array[17417] = 32'hFFFFFFF0;
    // rom_array[17418] = 32'hFFFFFFF0;
    // rom_array[17419] = 32'hFFFFFFF0;
    // rom_array[17420] = 32'hFFFFFFF0;
    // rom_array[17421] = 32'hFFFFFFF1;
    // rom_array[17422] = 32'hFFFFFFF1;
    // rom_array[17423] = 32'hFFFFFFF1;
    // rom_array[17424] = 32'hFFFFFFF1;
    // rom_array[17425] = 32'hFFFFFFF0;
    // rom_array[17426] = 32'hFFFFFFF0;
    // rom_array[17427] = 32'hFFFFFFF0;
    // rom_array[17428] = 32'hFFFFFFF0;
    // rom_array[17429] = 32'hFFFFFFF1;
    // rom_array[17430] = 32'hFFFFFFF1;
    // rom_array[17431] = 32'hFFFFFFF1;
    // rom_array[17432] = 32'hFFFFFFF1;
    // rom_array[17433] = 32'hFFFFFFF0;
    // rom_array[17434] = 32'hFFFFFFF0;
    // rom_array[17435] = 32'hFFFFFFF0;
    // rom_array[17436] = 32'hFFFFFFF0;
    // rom_array[17437] = 32'hFFFFFFF1;
    // rom_array[17438] = 32'hFFFFFFF1;
    // rom_array[17439] = 32'hFFFFFFF1;
    // rom_array[17440] = 32'hFFFFFFF1;
    // rom_array[17441] = 32'hFFFFFFF0;
    // rom_array[17442] = 32'hFFFFFFF0;
    // rom_array[17443] = 32'hFFFFFFF0;
    // rom_array[17444] = 32'hFFFFFFF0;
    // rom_array[17445] = 32'hFFFFFFF1;
    // rom_array[17446] = 32'hFFFFFFF1;
    // rom_array[17447] = 32'hFFFFFFF1;
    // rom_array[17448] = 32'hFFFFFFF1;
    // rom_array[17449] = 32'hFFFFFFF0;
    // rom_array[17450] = 32'hFFFFFFF0;
    // rom_array[17451] = 32'hFFFFFFF0;
    // rom_array[17452] = 32'hFFFFFFF0;
    // rom_array[17453] = 32'hFFFFFFF1;
    // rom_array[17454] = 32'hFFFFFFF1;
    // rom_array[17455] = 32'hFFFFFFF1;
    // rom_array[17456] = 32'hFFFFFFF1;
    // rom_array[17457] = 32'hFFFFFFF0;
    // rom_array[17458] = 32'hFFFFFFF0;
    // rom_array[17459] = 32'hFFFFFFF0;
    // rom_array[17460] = 32'hFFFFFFF0;
    // rom_array[17461] = 32'hFFFFFFF1;
    // rom_array[17462] = 32'hFFFFFFF1;
    // rom_array[17463] = 32'hFFFFFFF1;
    // rom_array[17464] = 32'hFFFFFFF1;
    // rom_array[17465] = 32'hFFFFFFF0;
    // rom_array[17466] = 32'hFFFFFFF0;
    // rom_array[17467] = 32'hFFFFFFF0;
    // rom_array[17468] = 32'hFFFFFFF0;
    // rom_array[17469] = 32'hFFFFFFF1;
    // rom_array[17470] = 32'hFFFFFFF1;
    // rom_array[17471] = 32'hFFFFFFF1;
    // rom_array[17472] = 32'hFFFFFFF1;
    // rom_array[17473] = 32'hFFFFFFF0;
    // rom_array[17474] = 32'hFFFFFFF0;
    // rom_array[17475] = 32'hFFFFFFF0;
    // rom_array[17476] = 32'hFFFFFFF0;
    // rom_array[17477] = 32'hFFFFFFF1;
    // rom_array[17478] = 32'hFFFFFFF1;
    // rom_array[17479] = 32'hFFFFFFF1;
    // rom_array[17480] = 32'hFFFFFFF1;
    // rom_array[17481] = 32'hFFFFFFF0;
    // rom_array[17482] = 32'hFFFFFFF0;
    // rom_array[17483] = 32'hFFFFFFF0;
    // rom_array[17484] = 32'hFFFFFFF0;
    // rom_array[17485] = 32'hFFFFFFF1;
    // rom_array[17486] = 32'hFFFFFFF1;
    // rom_array[17487] = 32'hFFFFFFF1;
    // rom_array[17488] = 32'hFFFFFFF1;
    // rom_array[17489] = 32'hFFFFFFF0;
    // rom_array[17490] = 32'hFFFFFFF0;
    // rom_array[17491] = 32'hFFFFFFF0;
    // rom_array[17492] = 32'hFFFFFFF0;
    // rom_array[17493] = 32'hFFFFFFF1;
    // rom_array[17494] = 32'hFFFFFFF1;
    // rom_array[17495] = 32'hFFFFFFF1;
    // rom_array[17496] = 32'hFFFFFFF1;
    // rom_array[17497] = 32'hFFFFFFF1;
    // rom_array[17498] = 32'hFFFFFFF1;
    // rom_array[17499] = 32'hFFFFFFF1;
    // rom_array[17500] = 32'hFFFFFFF1;
    // rom_array[17501] = 32'hFFFFFFF1;
    // rom_array[17502] = 32'hFFFFFFF1;
    // rom_array[17503] = 32'hFFFFFFF1;
    // rom_array[17504] = 32'hFFFFFFF1;
    // rom_array[17505] = 32'hFFFFFFF1;
    // rom_array[17506] = 32'hFFFFFFF1;
    // rom_array[17507] = 32'hFFFFFFF1;
    // rom_array[17508] = 32'hFFFFFFF1;
    // rom_array[17509] = 32'hFFFFFFF1;
    // rom_array[17510] = 32'hFFFFFFF1;
    // rom_array[17511] = 32'hFFFFFFF1;
    // rom_array[17512] = 32'hFFFFFFF1;
    // rom_array[17513] = 32'hFFFFFFF1;
    // rom_array[17514] = 32'hFFFFFFF1;
    // rom_array[17515] = 32'hFFFFFFF1;
    // rom_array[17516] = 32'hFFFFFFF1;
    // rom_array[17517] = 32'hFFFFFFF1;
    // rom_array[17518] = 32'hFFFFFFF1;
    // rom_array[17519] = 32'hFFFFFFF1;
    // rom_array[17520] = 32'hFFFFFFF1;
    // rom_array[17521] = 32'hFFFFFFF1;
    // rom_array[17522] = 32'hFFFFFFF1;
    // rom_array[17523] = 32'hFFFFFFF1;
    // rom_array[17524] = 32'hFFFFFFF1;
    // rom_array[17525] = 32'hFFFFFFF1;
    // rom_array[17526] = 32'hFFFFFFF1;
    // rom_array[17527] = 32'hFFFFFFF1;
    // rom_array[17528] = 32'hFFFFFFF1;
    // rom_array[17529] = 32'hFFFFFFF1;
    // rom_array[17530] = 32'hFFFFFFF1;
    // rom_array[17531] = 32'hFFFFFFF1;
    // rom_array[17532] = 32'hFFFFFFF1;
    // rom_array[17533] = 32'hFFFFFFF1;
    // rom_array[17534] = 32'hFFFFFFF1;
    // rom_array[17535] = 32'hFFFFFFF1;
    // rom_array[17536] = 32'hFFFFFFF1;
    // rom_array[17537] = 32'hFFFFFFF1;
    // rom_array[17538] = 32'hFFFFFFF1;
    // rom_array[17539] = 32'hFFFFFFF1;
    // rom_array[17540] = 32'hFFFFFFF1;
    // rom_array[17541] = 32'hFFFFFFF1;
    // rom_array[17542] = 32'hFFFFFFF1;
    // rom_array[17543] = 32'hFFFFFFF1;
    // rom_array[17544] = 32'hFFFFFFF1;
    // rom_array[17545] = 32'hFFFFFFF1;
    // rom_array[17546] = 32'hFFFFFFF1;
    // rom_array[17547] = 32'hFFFFFFF1;
    // rom_array[17548] = 32'hFFFFFFF1;
    // rom_array[17549] = 32'hFFFFFFF0;
    // rom_array[17550] = 32'hFFFFFFF0;
    // rom_array[17551] = 32'hFFFFFFF0;
    // rom_array[17552] = 32'hFFFFFFF0;
    // rom_array[17553] = 32'hFFFFFFF1;
    // rom_array[17554] = 32'hFFFFFFF1;
    // rom_array[17555] = 32'hFFFFFFF1;
    // rom_array[17556] = 32'hFFFFFFF1;
    // rom_array[17557] = 32'hFFFFFFF0;
    // rom_array[17558] = 32'hFFFFFFF0;
    // rom_array[17559] = 32'hFFFFFFF0;
    // rom_array[17560] = 32'hFFFFFFF0;
    // rom_array[17561] = 32'hFFFFFFF1;
    // rom_array[17562] = 32'hFFFFFFF1;
    // rom_array[17563] = 32'hFFFFFFF1;
    // rom_array[17564] = 32'hFFFFFFF1;
    // rom_array[17565] = 32'hFFFFFFF1;
    // rom_array[17566] = 32'hFFFFFFF1;
    // rom_array[17567] = 32'hFFFFFFF1;
    // rom_array[17568] = 32'hFFFFFFF1;
    // rom_array[17569] = 32'hFFFFFFF1;
    // rom_array[17570] = 32'hFFFFFFF1;
    // rom_array[17571] = 32'hFFFFFFF1;
    // rom_array[17572] = 32'hFFFFFFF1;
    // rom_array[17573] = 32'hFFFFFFF1;
    // rom_array[17574] = 32'hFFFFFFF1;
    // rom_array[17575] = 32'hFFFFFFF1;
    // rom_array[17576] = 32'hFFFFFFF1;
    // rom_array[17577] = 32'hFFFFFFF1;
    // rom_array[17578] = 32'hFFFFFFF1;
    // rom_array[17579] = 32'hFFFFFFF1;
    // rom_array[17580] = 32'hFFFFFFF1;
    // rom_array[17581] = 32'hFFFFFFF0;
    // rom_array[17582] = 32'hFFFFFFF0;
    // rom_array[17583] = 32'hFFFFFFF0;
    // rom_array[17584] = 32'hFFFFFFF0;
    // rom_array[17585] = 32'hFFFFFFF1;
    // rom_array[17586] = 32'hFFFFFFF1;
    // rom_array[17587] = 32'hFFFFFFF1;
    // rom_array[17588] = 32'hFFFFFFF1;
    // rom_array[17589] = 32'hFFFFFFF0;
    // rom_array[17590] = 32'hFFFFFFF0;
    // rom_array[17591] = 32'hFFFFFFF0;
    // rom_array[17592] = 32'hFFFFFFF0;
    // rom_array[17593] = 32'hFFFFFFF1;
    // rom_array[17594] = 32'hFFFFFFF1;
    // rom_array[17595] = 32'hFFFFFFF1;
    // rom_array[17596] = 32'hFFFFFFF1;
    // rom_array[17597] = 32'hFFFFFFF0;
    // rom_array[17598] = 32'hFFFFFFF0;
    // rom_array[17599] = 32'hFFFFFFF0;
    // rom_array[17600] = 32'hFFFFFFF0;
    // rom_array[17601] = 32'hFFFFFFF1;
    // rom_array[17602] = 32'hFFFFFFF1;
    // rom_array[17603] = 32'hFFFFFFF1;
    // rom_array[17604] = 32'hFFFFFFF1;
    // rom_array[17605] = 32'hFFFFFFF0;
    // rom_array[17606] = 32'hFFFFFFF0;
    // rom_array[17607] = 32'hFFFFFFF0;
    // rom_array[17608] = 32'hFFFFFFF0;
    // rom_array[17609] = 32'hFFFFFFF1;
    // rom_array[17610] = 32'hFFFFFFF1;
    // rom_array[17611] = 32'hFFFFFFF1;
    // rom_array[17612] = 32'hFFFFFFF1;
    // rom_array[17613] = 32'hFFFFFFF0;
    // rom_array[17614] = 32'hFFFFFFF0;
    // rom_array[17615] = 32'hFFFFFFF0;
    // rom_array[17616] = 32'hFFFFFFF0;
    // rom_array[17617] = 32'hFFFFFFF1;
    // rom_array[17618] = 32'hFFFFFFF1;
    // rom_array[17619] = 32'hFFFFFFF1;
    // rom_array[17620] = 32'hFFFFFFF1;
    // rom_array[17621] = 32'hFFFFFFF0;
    // rom_array[17622] = 32'hFFFFFFF0;
    // rom_array[17623] = 32'hFFFFFFF0;
    // rom_array[17624] = 32'hFFFFFFF0;
    // rom_array[17625] = 32'hFFFFFFF1;
    // rom_array[17626] = 32'hFFFFFFF1;
    // rom_array[17627] = 32'hFFFFFFF1;
    // rom_array[17628] = 32'hFFFFFFF1;
    // rom_array[17629] = 32'hFFFFFFF0;
    // rom_array[17630] = 32'hFFFFFFF0;
    // rom_array[17631] = 32'hFFFFFFF0;
    // rom_array[17632] = 32'hFFFFFFF0;
    // rom_array[17633] = 32'hFFFFFFF1;
    // rom_array[17634] = 32'hFFFFFFF1;
    // rom_array[17635] = 32'hFFFFFFF1;
    // rom_array[17636] = 32'hFFFFFFF1;
    // rom_array[17637] = 32'hFFFFFFF0;
    // rom_array[17638] = 32'hFFFFFFF0;
    // rom_array[17639] = 32'hFFFFFFF0;
    // rom_array[17640] = 32'hFFFFFFF0;
    // rom_array[17641] = 32'hFFFFFFF1;
    // rom_array[17642] = 32'hFFFFFFF1;
    // rom_array[17643] = 32'hFFFFFFF1;
    // rom_array[17644] = 32'hFFFFFFF1;
    // rom_array[17645] = 32'hFFFFFFF0;
    // rom_array[17646] = 32'hFFFFFFF0;
    // rom_array[17647] = 32'hFFFFFFF0;
    // rom_array[17648] = 32'hFFFFFFF0;
    // rom_array[17649] = 32'hFFFFFFF1;
    // rom_array[17650] = 32'hFFFFFFF1;
    // rom_array[17651] = 32'hFFFFFFF1;
    // rom_array[17652] = 32'hFFFFFFF1;
    // rom_array[17653] = 32'hFFFFFFF0;
    // rom_array[17654] = 32'hFFFFFFF0;
    // rom_array[17655] = 32'hFFFFFFF0;
    // rom_array[17656] = 32'hFFFFFFF0;
    // rom_array[17657] = 32'hFFFFFFF1;
    // rom_array[17658] = 32'hFFFFFFF1;
    // rom_array[17659] = 32'hFFFFFFF1;
    // rom_array[17660] = 32'hFFFFFFF1;
    // rom_array[17661] = 32'hFFFFFFF0;
    // rom_array[17662] = 32'hFFFFFFF0;
    // rom_array[17663] = 32'hFFFFFFF0;
    // rom_array[17664] = 32'hFFFFFFF0;
    // rom_array[17665] = 32'hFFFFFFF1;
    // rom_array[17666] = 32'hFFFFFFF1;
    // rom_array[17667] = 32'hFFFFFFF1;
    // rom_array[17668] = 32'hFFFFFFF1;
    // rom_array[17669] = 32'hFFFFFFF0;
    // rom_array[17670] = 32'hFFFFFFF0;
    // rom_array[17671] = 32'hFFFFFFF0;
    // rom_array[17672] = 32'hFFFFFFF0;
    // rom_array[17673] = 32'hFFFFFFF0;
    // rom_array[17674] = 32'hFFFFFFF0;
    // rom_array[17675] = 32'hFFFFFFF1;
    // rom_array[17676] = 32'hFFFFFFF1;
    // rom_array[17677] = 32'hFFFFFFF0;
    // rom_array[17678] = 32'hFFFFFFF0;
    // rom_array[17679] = 32'hFFFFFFF1;
    // rom_array[17680] = 32'hFFFFFFF1;
    // rom_array[17681] = 32'hFFFFFFF0;
    // rom_array[17682] = 32'hFFFFFFF0;
    // rom_array[17683] = 32'hFFFFFFF1;
    // rom_array[17684] = 32'hFFFFFFF1;
    // rom_array[17685] = 32'hFFFFFFF0;
    // rom_array[17686] = 32'hFFFFFFF0;
    // rom_array[17687] = 32'hFFFFFFF1;
    // rom_array[17688] = 32'hFFFFFFF1;
    // rom_array[17689] = 32'hFFFFFFF0;
    // rom_array[17690] = 32'hFFFFFFF0;
    // rom_array[17691] = 32'hFFFFFFF1;
    // rom_array[17692] = 32'hFFFFFFF1;
    // rom_array[17693] = 32'hFFFFFFF0;
    // rom_array[17694] = 32'hFFFFFFF0;
    // rom_array[17695] = 32'hFFFFFFF1;
    // rom_array[17696] = 32'hFFFFFFF1;
    // rom_array[17697] = 32'hFFFFFFF0;
    // rom_array[17698] = 32'hFFFFFFF0;
    // rom_array[17699] = 32'hFFFFFFF1;
    // rom_array[17700] = 32'hFFFFFFF1;
    // rom_array[17701] = 32'hFFFFFFF0;
    // rom_array[17702] = 32'hFFFFFFF0;
    // rom_array[17703] = 32'hFFFFFFF1;
    // rom_array[17704] = 32'hFFFFFFF1;
    // rom_array[17705] = 32'hFFFFFFF0;
    // rom_array[17706] = 32'hFFFFFFF0;
    // rom_array[17707] = 32'hFFFFFFF1;
    // rom_array[17708] = 32'hFFFFFFF1;
    // rom_array[17709] = 32'hFFFFFFF0;
    // rom_array[17710] = 32'hFFFFFFF0;
    // rom_array[17711] = 32'hFFFFFFF1;
    // rom_array[17712] = 32'hFFFFFFF1;
    // rom_array[17713] = 32'hFFFFFFF0;
    // rom_array[17714] = 32'hFFFFFFF0;
    // rom_array[17715] = 32'hFFFFFFF1;
    // rom_array[17716] = 32'hFFFFFFF1;
    // rom_array[17717] = 32'hFFFFFFF0;
    // rom_array[17718] = 32'hFFFFFFF0;
    // rom_array[17719] = 32'hFFFFFFF1;
    // rom_array[17720] = 32'hFFFFFFF1;
    // rom_array[17721] = 32'hFFFFFFF0;
    // rom_array[17722] = 32'hFFFFFFF0;
    // rom_array[17723] = 32'hFFFFFFF1;
    // rom_array[17724] = 32'hFFFFFFF1;
    // rom_array[17725] = 32'hFFFFFFF0;
    // rom_array[17726] = 32'hFFFFFFF0;
    // rom_array[17727] = 32'hFFFFFFF0;
    // rom_array[17728] = 32'hFFFFFFF0;
    // rom_array[17729] = 32'hFFFFFFF0;
    // rom_array[17730] = 32'hFFFFFFF0;
    // rom_array[17731] = 32'hFFFFFFF1;
    // rom_array[17732] = 32'hFFFFFFF1;
    // rom_array[17733] = 32'hFFFFFFF0;
    // rom_array[17734] = 32'hFFFFFFF0;
    // rom_array[17735] = 32'hFFFFFFF0;
    // rom_array[17736] = 32'hFFFFFFF0;
    // rom_array[17737] = 32'hFFFFFFF1;
    // rom_array[17738] = 32'hFFFFFFF1;
    // rom_array[17739] = 32'hFFFFFFF1;
    // rom_array[17740] = 32'hFFFFFFF1;
    // rom_array[17741] = 32'hFFFFFFF0;
    // rom_array[17742] = 32'hFFFFFFF0;
    // rom_array[17743] = 32'hFFFFFFF0;
    // rom_array[17744] = 32'hFFFFFFF0;
    // rom_array[17745] = 32'hFFFFFFF1;
    // rom_array[17746] = 32'hFFFFFFF1;
    // rom_array[17747] = 32'hFFFFFFF1;
    // rom_array[17748] = 32'hFFFFFFF1;
    // rom_array[17749] = 32'hFFFFFFF0;
    // rom_array[17750] = 32'hFFFFFFF0;
    // rom_array[17751] = 32'hFFFFFFF0;
    // rom_array[17752] = 32'hFFFFFFF0;
    // rom_array[17753] = 32'hFFFFFFF1;
    // rom_array[17754] = 32'hFFFFFFF1;
    // rom_array[17755] = 32'hFFFFFFF1;
    // rom_array[17756] = 32'hFFFFFFF1;
    // rom_array[17757] = 32'hFFFFFFF0;
    // rom_array[17758] = 32'hFFFFFFF0;
    // rom_array[17759] = 32'hFFFFFFF0;
    // rom_array[17760] = 32'hFFFFFFF0;
    // rom_array[17761] = 32'hFFFFFFF1;
    // rom_array[17762] = 32'hFFFFFFF1;
    // rom_array[17763] = 32'hFFFFFFF1;
    // rom_array[17764] = 32'hFFFFFFF1;
    // rom_array[17765] = 32'hFFFFFFF0;
    // rom_array[17766] = 32'hFFFFFFF0;
    // rom_array[17767] = 32'hFFFFFFF0;
    // rom_array[17768] = 32'hFFFFFFF0;
    // rom_array[17769] = 32'hFFFFFFF1;
    // rom_array[17770] = 32'hFFFFFFF1;
    // rom_array[17771] = 32'hFFFFFFF1;
    // rom_array[17772] = 32'hFFFFFFF1;
    // rom_array[17773] = 32'hFFFFFFF0;
    // rom_array[17774] = 32'hFFFFFFF0;
    // rom_array[17775] = 32'hFFFFFFF0;
    // rom_array[17776] = 32'hFFFFFFF0;
    // rom_array[17777] = 32'hFFFFFFF1;
    // rom_array[17778] = 32'hFFFFFFF1;
    // rom_array[17779] = 32'hFFFFFFF1;
    // rom_array[17780] = 32'hFFFFFFF1;
    // rom_array[17781] = 32'hFFFFFFF0;
    // rom_array[17782] = 32'hFFFFFFF0;
    // rom_array[17783] = 32'hFFFFFFF0;
    // rom_array[17784] = 32'hFFFFFFF0;
    // rom_array[17785] = 32'hFFFFFFF1;
    // rom_array[17786] = 32'hFFFFFFF1;
    // rom_array[17787] = 32'hFFFFFFF1;
    // rom_array[17788] = 32'hFFFFFFF1;
    // rom_array[17789] = 32'hFFFFFFF1;
    // rom_array[17790] = 32'hFFFFFFF1;
    // rom_array[17791] = 32'hFFFFFFF1;
    // rom_array[17792] = 32'hFFFFFFF1;
    // rom_array[17793] = 32'hFFFFFFF1;
    // rom_array[17794] = 32'hFFFFFFF1;
    // rom_array[17795] = 32'hFFFFFFF1;
    // rom_array[17796] = 32'hFFFFFFF1;
    // rom_array[17797] = 32'hFFFFFFF1;
    // rom_array[17798] = 32'hFFFFFFF1;
    // rom_array[17799] = 32'hFFFFFFF1;
    // rom_array[17800] = 32'hFFFFFFF1;
    // rom_array[17801] = 32'hFFFFFFF1;
    // rom_array[17802] = 32'hFFFFFFF1;
    // rom_array[17803] = 32'hFFFFFFF1;
    // rom_array[17804] = 32'hFFFFFFF1;
    // rom_array[17805] = 32'hFFFFFFF1;
    // rom_array[17806] = 32'hFFFFFFF1;
    // rom_array[17807] = 32'hFFFFFFF1;
    // rom_array[17808] = 32'hFFFFFFF1;
    // rom_array[17809] = 32'hFFFFFFF1;
    // rom_array[17810] = 32'hFFFFFFF1;
    // rom_array[17811] = 32'hFFFFFFF1;
    // rom_array[17812] = 32'hFFFFFFF1;
    // rom_array[17813] = 32'hFFFFFFF1;
    // rom_array[17814] = 32'hFFFFFFF1;
    // rom_array[17815] = 32'hFFFFFFF1;
    // rom_array[17816] = 32'hFFFFFFF1;
    // rom_array[17817] = 32'hFFFFFFF1;
    // rom_array[17818] = 32'hFFFFFFF1;
    // rom_array[17819] = 32'hFFFFFFF1;
    // rom_array[17820] = 32'hFFFFFFF1;
    // rom_array[17821] = 32'hFFFFFFF1;
    // rom_array[17822] = 32'hFFFFFFF1;
    // rom_array[17823] = 32'hFFFFFFF1;
    // rom_array[17824] = 32'hFFFFFFF1;
    // rom_array[17825] = 32'hFFFFFFF1;
    // rom_array[17826] = 32'hFFFFFFF1;
    // rom_array[17827] = 32'hFFFFFFF1;
    // rom_array[17828] = 32'hFFFFFFF1;
    // rom_array[17829] = 32'hFFFFFFF1;
    // rom_array[17830] = 32'hFFFFFFF1;
    // rom_array[17831] = 32'hFFFFFFF1;
    // rom_array[17832] = 32'hFFFFFFF1;
    // rom_array[17833] = 32'hFFFFFFF1;
    // rom_array[17834] = 32'hFFFFFFF1;
    // rom_array[17835] = 32'hFFFFFFF1;
    // rom_array[17836] = 32'hFFFFFFF1;
    // rom_array[17837] = 32'hFFFFFFF0;
    // rom_array[17838] = 32'hFFFFFFF0;
    // rom_array[17839] = 32'hFFFFFFF0;
    // rom_array[17840] = 32'hFFFFFFF0;
    // rom_array[17841] = 32'hFFFFFFF1;
    // rom_array[17842] = 32'hFFFFFFF1;
    // rom_array[17843] = 32'hFFFFFFF1;
    // rom_array[17844] = 32'hFFFFFFF1;
    // rom_array[17845] = 32'hFFFFFFF0;
    // rom_array[17846] = 32'hFFFFFFF0;
    // rom_array[17847] = 32'hFFFFFFF0;
    // rom_array[17848] = 32'hFFFFFFF0;
    // rom_array[17849] = 32'hFFFFFFF0;
    // rom_array[17850] = 32'hFFFFFFF0;
    // rom_array[17851] = 32'hFFFFFFF0;
    // rom_array[17852] = 32'hFFFFFFF0;
    // rom_array[17853] = 32'hFFFFFFF0;
    // rom_array[17854] = 32'hFFFFFFF0;
    // rom_array[17855] = 32'hFFFFFFF1;
    // rom_array[17856] = 32'hFFFFFFF1;
    // rom_array[17857] = 32'hFFFFFFF0;
    // rom_array[17858] = 32'hFFFFFFF0;
    // rom_array[17859] = 32'hFFFFFFF0;
    // rom_array[17860] = 32'hFFFFFFF0;
    // rom_array[17861] = 32'hFFFFFFF0;
    // rom_array[17862] = 32'hFFFFFFF0;
    // rom_array[17863] = 32'hFFFFFFF1;
    // rom_array[17864] = 32'hFFFFFFF1;
    // rom_array[17865] = 32'hFFFFFFF0;
    // rom_array[17866] = 32'hFFFFFFF0;
    // rom_array[17867] = 32'hFFFFFFF0;
    // rom_array[17868] = 32'hFFFFFFF0;
    // rom_array[17869] = 32'hFFFFFFF1;
    // rom_array[17870] = 32'hFFFFFFF1;
    // rom_array[17871] = 32'hFFFFFFF1;
    // rom_array[17872] = 32'hFFFFFFF1;
    // rom_array[17873] = 32'hFFFFFFF0;
    // rom_array[17874] = 32'hFFFFFFF0;
    // rom_array[17875] = 32'hFFFFFFF0;
    // rom_array[17876] = 32'hFFFFFFF0;
    // rom_array[17877] = 32'hFFFFFFF1;
    // rom_array[17878] = 32'hFFFFFFF1;
    // rom_array[17879] = 32'hFFFFFFF1;
    // rom_array[17880] = 32'hFFFFFFF1;
    // rom_array[17881] = 32'hFFFFFFF0;
    // rom_array[17882] = 32'hFFFFFFF0;
    // rom_array[17883] = 32'hFFFFFFF1;
    // rom_array[17884] = 32'hFFFFFFF1;
    // rom_array[17885] = 32'hFFFFFFF0;
    // rom_array[17886] = 32'hFFFFFFF0;
    // rom_array[17887] = 32'hFFFFFFF1;
    // rom_array[17888] = 32'hFFFFFFF1;
    // rom_array[17889] = 32'hFFFFFFF0;
    // rom_array[17890] = 32'hFFFFFFF0;
    // rom_array[17891] = 32'hFFFFFFF1;
    // rom_array[17892] = 32'hFFFFFFF1;
    // rom_array[17893] = 32'hFFFFFFF0;
    // rom_array[17894] = 32'hFFFFFFF0;
    // rom_array[17895] = 32'hFFFFFFF1;
    // rom_array[17896] = 32'hFFFFFFF1;
    // rom_array[17897] = 32'hFFFFFFF0;
    // rom_array[17898] = 32'hFFFFFFF0;
    // rom_array[17899] = 32'hFFFFFFF0;
    // rom_array[17900] = 32'hFFFFFFF0;
    // rom_array[17901] = 32'hFFFFFFF1;
    // rom_array[17902] = 32'hFFFFFFF1;
    // rom_array[17903] = 32'hFFFFFFF1;
    // rom_array[17904] = 32'hFFFFFFF1;
    // rom_array[17905] = 32'hFFFFFFF0;
    // rom_array[17906] = 32'hFFFFFFF0;
    // rom_array[17907] = 32'hFFFFFFF0;
    // rom_array[17908] = 32'hFFFFFFF0;
    // rom_array[17909] = 32'hFFFFFFF1;
    // rom_array[17910] = 32'hFFFFFFF1;
    // rom_array[17911] = 32'hFFFFFFF1;
    // rom_array[17912] = 32'hFFFFFFF1;
    // rom_array[17913] = 32'hFFFFFFF0;
    // rom_array[17914] = 32'hFFFFFFF0;
    // rom_array[17915] = 32'hFFFFFFF0;
    // rom_array[17916] = 32'hFFFFFFF0;
    // rom_array[17917] = 32'hFFFFFFF1;
    // rom_array[17918] = 32'hFFFFFFF1;
    // rom_array[17919] = 32'hFFFFFFF1;
    // rom_array[17920] = 32'hFFFFFFF1;
    // rom_array[17921] = 32'hFFFFFFF0;
    // rom_array[17922] = 32'hFFFFFFF0;
    // rom_array[17923] = 32'hFFFFFFF0;
    // rom_array[17924] = 32'hFFFFFFF0;
    // rom_array[17925] = 32'hFFFFFFF1;
    // rom_array[17926] = 32'hFFFFFFF1;
    // rom_array[17927] = 32'hFFFFFFF1;
    // rom_array[17928] = 32'hFFFFFFF1;
    // rom_array[17929] = 32'hFFFFFFF0;
    // rom_array[17930] = 32'hFFFFFFF0;
    // rom_array[17931] = 32'hFFFFFFF0;
    // rom_array[17932] = 32'hFFFFFFF0;
    // rom_array[17933] = 32'hFFFFFFF1;
    // rom_array[17934] = 32'hFFFFFFF1;
    // rom_array[17935] = 32'hFFFFFFF1;
    // rom_array[17936] = 32'hFFFFFFF1;
    // rom_array[17937] = 32'hFFFFFFF0;
    // rom_array[17938] = 32'hFFFFFFF0;
    // rom_array[17939] = 32'hFFFFFFF0;
    // rom_array[17940] = 32'hFFFFFFF0;
    // rom_array[17941] = 32'hFFFFFFF1;
    // rom_array[17942] = 32'hFFFFFFF1;
    // rom_array[17943] = 32'hFFFFFFF1;
    // rom_array[17944] = 32'hFFFFFFF1;
    // rom_array[17945] = 32'hFFFFFFF0;
    // rom_array[17946] = 32'hFFFFFFF0;
    // rom_array[17947] = 32'hFFFFFFF0;
    // rom_array[17948] = 32'hFFFFFFF0;
    // rom_array[17949] = 32'hFFFFFFF1;
    // rom_array[17950] = 32'hFFFFFFF1;
    // rom_array[17951] = 32'hFFFFFFF1;
    // rom_array[17952] = 32'hFFFFFFF1;
    // rom_array[17953] = 32'hFFFFFFF0;
    // rom_array[17954] = 32'hFFFFFFF0;
    // rom_array[17955] = 32'hFFFFFFF0;
    // rom_array[17956] = 32'hFFFFFFF0;
    // rom_array[17957] = 32'hFFFFFFF1;
    // rom_array[17958] = 32'hFFFFFFF1;
    // rom_array[17959] = 32'hFFFFFFF1;
    // rom_array[17960] = 32'hFFFFFFF1;
    // rom_array[17961] = 32'hFFFFFFF0;
    // rom_array[17962] = 32'hFFFFFFF0;
    // rom_array[17963] = 32'hFFFFFFF0;
    // rom_array[17964] = 32'hFFFFFFF0;
    // rom_array[17965] = 32'hFFFFFFF1;
    // rom_array[17966] = 32'hFFFFFFF1;
    // rom_array[17967] = 32'hFFFFFFF1;
    // rom_array[17968] = 32'hFFFFFFF1;
    // rom_array[17969] = 32'hFFFFFFF0;
    // rom_array[17970] = 32'hFFFFFFF0;
    // rom_array[17971] = 32'hFFFFFFF0;
    // rom_array[17972] = 32'hFFFFFFF0;
    // rom_array[17973] = 32'hFFFFFFF1;
    // rom_array[17974] = 32'hFFFFFFF1;
    // rom_array[17975] = 32'hFFFFFFF1;
    // rom_array[17976] = 32'hFFFFFFF1;
    // rom_array[17977] = 32'hFFFFFFF0;
    // rom_array[17978] = 32'hFFFFFFF0;
    // rom_array[17979] = 32'hFFFFFFF0;
    // rom_array[17980] = 32'hFFFFFFF0;
    // rom_array[17981] = 32'hFFFFFFF1;
    // rom_array[17982] = 32'hFFFFFFF1;
    // rom_array[17983] = 32'hFFFFFFF1;
    // rom_array[17984] = 32'hFFFFFFF1;
    // rom_array[17985] = 32'hFFFFFFF0;
    // rom_array[17986] = 32'hFFFFFFF0;
    // rom_array[17987] = 32'hFFFFFFF0;
    // rom_array[17988] = 32'hFFFFFFF0;
    // rom_array[17989] = 32'hFFFFFFF1;
    // rom_array[17990] = 32'hFFFFFFF1;
    // rom_array[17991] = 32'hFFFFFFF1;
    // rom_array[17992] = 32'hFFFFFFF1;
    // rom_array[17993] = 32'hFFFFFFF1;
    // rom_array[17994] = 32'hFFFFFFF1;
    // rom_array[17995] = 32'hFFFFFFF1;
    // rom_array[17996] = 32'hFFFFFFF1;
    // rom_array[17997] = 32'hFFFFFFF1;
    // rom_array[17998] = 32'hFFFFFFF1;
    // rom_array[17999] = 32'hFFFFFFF1;
    // rom_array[18000] = 32'hFFFFFFF1;
    // rom_array[18001] = 32'hFFFFFFF1;
    // rom_array[18002] = 32'hFFFFFFF1;
    // rom_array[18003] = 32'hFFFFFFF1;
    // rom_array[18004] = 32'hFFFFFFF1;
    // rom_array[18005] = 32'hFFFFFFF1;
    // rom_array[18006] = 32'hFFFFFFF1;
    // rom_array[18007] = 32'hFFFFFFF1;
    // rom_array[18008] = 32'hFFFFFFF1;
    // rom_array[18009] = 32'hFFFFFFF0;
    // rom_array[18010] = 32'hFFFFFFF0;
    // rom_array[18011] = 32'hFFFFFFF0;
    // rom_array[18012] = 32'hFFFFFFF0;
    // rom_array[18013] = 32'hFFFFFFF1;
    // rom_array[18014] = 32'hFFFFFFF1;
    // rom_array[18015] = 32'hFFFFFFF1;
    // rom_array[18016] = 32'hFFFFFFF1;
    // rom_array[18017] = 32'hFFFFFFF0;
    // rom_array[18018] = 32'hFFFFFFF0;
    // rom_array[18019] = 32'hFFFFFFF0;
    // rom_array[18020] = 32'hFFFFFFF0;
    // rom_array[18021] = 32'hFFFFFFF1;
    // rom_array[18022] = 32'hFFFFFFF1;
    // rom_array[18023] = 32'hFFFFFFF1;
    // rom_array[18024] = 32'hFFFFFFF1;
    // rom_array[18025] = 32'hFFFFFFF0;
    // rom_array[18026] = 32'hFFFFFFF0;
    // rom_array[18027] = 32'hFFFFFFF0;
    // rom_array[18028] = 32'hFFFFFFF0;
    // rom_array[18029] = 32'hFFFFFFF1;
    // rom_array[18030] = 32'hFFFFFFF1;
    // rom_array[18031] = 32'hFFFFFFF1;
    // rom_array[18032] = 32'hFFFFFFF1;
    // rom_array[18033] = 32'hFFFFFFF0;
    // rom_array[18034] = 32'hFFFFFFF0;
    // rom_array[18035] = 32'hFFFFFFF0;
    // rom_array[18036] = 32'hFFFFFFF0;
    // rom_array[18037] = 32'hFFFFFFF1;
    // rom_array[18038] = 32'hFFFFFFF1;
    // rom_array[18039] = 32'hFFFFFFF1;
    // rom_array[18040] = 32'hFFFFFFF1;
    // rom_array[18041] = 32'hFFFFFFF1;
    // rom_array[18042] = 32'hFFFFFFF1;
    // rom_array[18043] = 32'hFFFFFFF1;
    // rom_array[18044] = 32'hFFFFFFF1;
    // rom_array[18045] = 32'hFFFFFFF1;
    // rom_array[18046] = 32'hFFFFFFF1;
    // rom_array[18047] = 32'hFFFFFFF1;
    // rom_array[18048] = 32'hFFFFFFF1;
    // rom_array[18049] = 32'hFFFFFFF1;
    // rom_array[18050] = 32'hFFFFFFF1;
    // rom_array[18051] = 32'hFFFFFFF1;
    // rom_array[18052] = 32'hFFFFFFF1;
    // rom_array[18053] = 32'hFFFFFFF1;
    // rom_array[18054] = 32'hFFFFFFF1;
    // rom_array[18055] = 32'hFFFFFFF1;
    // rom_array[18056] = 32'hFFFFFFF1;
    // rom_array[18057] = 32'hFFFFFFF1;
    // rom_array[18058] = 32'hFFFFFFF1;
    // rom_array[18059] = 32'hFFFFFFF1;
    // rom_array[18060] = 32'hFFFFFFF1;
    // rom_array[18061] = 32'hFFFFFFF1;
    // rom_array[18062] = 32'hFFFFFFF1;
    // rom_array[18063] = 32'hFFFFFFF1;
    // rom_array[18064] = 32'hFFFFFFF1;
    // rom_array[18065] = 32'hFFFFFFF1;
    // rom_array[18066] = 32'hFFFFFFF1;
    // rom_array[18067] = 32'hFFFFFFF1;
    // rom_array[18068] = 32'hFFFFFFF1;
    // rom_array[18069] = 32'hFFFFFFF1;
    // rom_array[18070] = 32'hFFFFFFF1;
    // rom_array[18071] = 32'hFFFFFFF1;
    // rom_array[18072] = 32'hFFFFFFF1;
    // rom_array[18073] = 32'hFFFFFFF0;
    // rom_array[18074] = 32'hFFFFFFF0;
    // rom_array[18075] = 32'hFFFFFFF0;
    // rom_array[18076] = 32'hFFFFFFF0;
    // rom_array[18077] = 32'hFFFFFFF1;
    // rom_array[18078] = 32'hFFFFFFF1;
    // rom_array[18079] = 32'hFFFFFFF1;
    // rom_array[18080] = 32'hFFFFFFF1;
    // rom_array[18081] = 32'hFFFFFFF0;
    // rom_array[18082] = 32'hFFFFFFF0;
    // rom_array[18083] = 32'hFFFFFFF0;
    // rom_array[18084] = 32'hFFFFFFF0;
    // rom_array[18085] = 32'hFFFFFFF1;
    // rom_array[18086] = 32'hFFFFFFF1;
    // rom_array[18087] = 32'hFFFFFFF1;
    // rom_array[18088] = 32'hFFFFFFF1;
    // rom_array[18089] = 32'hFFFFFFF0;
    // rom_array[18090] = 32'hFFFFFFF0;
    // rom_array[18091] = 32'hFFFFFFF0;
    // rom_array[18092] = 32'hFFFFFFF0;
    // rom_array[18093] = 32'hFFFFFFF1;
    // rom_array[18094] = 32'hFFFFFFF1;
    // rom_array[18095] = 32'hFFFFFFF1;
    // rom_array[18096] = 32'hFFFFFFF1;
    // rom_array[18097] = 32'hFFFFFFF0;
    // rom_array[18098] = 32'hFFFFFFF0;
    // rom_array[18099] = 32'hFFFFFFF0;
    // rom_array[18100] = 32'hFFFFFFF0;
    // rom_array[18101] = 32'hFFFFFFF1;
    // rom_array[18102] = 32'hFFFFFFF1;
    // rom_array[18103] = 32'hFFFFFFF1;
    // rom_array[18104] = 32'hFFFFFFF1;
    // rom_array[18105] = 32'hFFFFFFF1;
    // rom_array[18106] = 32'hFFFFFFF1;
    // rom_array[18107] = 32'hFFFFFFF1;
    // rom_array[18108] = 32'hFFFFFFF1;
    // rom_array[18109] = 32'hFFFFFFF1;
    // rom_array[18110] = 32'hFFFFFFF1;
    // rom_array[18111] = 32'hFFFFFFF1;
    // rom_array[18112] = 32'hFFFFFFF1;
    // rom_array[18113] = 32'hFFFFFFF1;
    // rom_array[18114] = 32'hFFFFFFF1;
    // rom_array[18115] = 32'hFFFFFFF1;
    // rom_array[18116] = 32'hFFFFFFF1;
    // rom_array[18117] = 32'hFFFFFFF1;
    // rom_array[18118] = 32'hFFFFFFF1;
    // rom_array[18119] = 32'hFFFFFFF1;
    // rom_array[18120] = 32'hFFFFFFF1;
    // rom_array[18121] = 32'hFFFFFFF1;
    // rom_array[18122] = 32'hFFFFFFF1;
    // rom_array[18123] = 32'hFFFFFFF1;
    // rom_array[18124] = 32'hFFFFFFF1;
    // rom_array[18125] = 32'hFFFFFFF1;
    // rom_array[18126] = 32'hFFFFFFF1;
    // rom_array[18127] = 32'hFFFFFFF1;
    // rom_array[18128] = 32'hFFFFFFF1;
    // rom_array[18129] = 32'hFFFFFFF1;
    // rom_array[18130] = 32'hFFFFFFF1;
    // rom_array[18131] = 32'hFFFFFFF1;
    // rom_array[18132] = 32'hFFFFFFF1;
    // rom_array[18133] = 32'hFFFFFFF1;
    // rom_array[18134] = 32'hFFFFFFF1;
    // rom_array[18135] = 32'hFFFFFFF1;
    // rom_array[18136] = 32'hFFFFFFF1;
    // rom_array[18137] = 32'hFFFFFFF0;
    // rom_array[18138] = 32'hFFFFFFF0;
    // rom_array[18139] = 32'hFFFFFFF1;
    // rom_array[18140] = 32'hFFFFFFF1;
    // rom_array[18141] = 32'hFFFFFFF0;
    // rom_array[18142] = 32'hFFFFFFF0;
    // rom_array[18143] = 32'hFFFFFFF1;
    // rom_array[18144] = 32'hFFFFFFF1;
    // rom_array[18145] = 32'hFFFFFFF0;
    // rom_array[18146] = 32'hFFFFFFF0;
    // rom_array[18147] = 32'hFFFFFFF1;
    // rom_array[18148] = 32'hFFFFFFF1;
    // rom_array[18149] = 32'hFFFFFFF0;
    // rom_array[18150] = 32'hFFFFFFF0;
    // rom_array[18151] = 32'hFFFFFFF1;
    // rom_array[18152] = 32'hFFFFFFF1;
    // rom_array[18153] = 32'hFFFFFFF0;
    // rom_array[18154] = 32'hFFFFFFF0;
    // rom_array[18155] = 32'hFFFFFFF1;
    // rom_array[18156] = 32'hFFFFFFF1;
    // rom_array[18157] = 32'hFFFFFFF0;
    // rom_array[18158] = 32'hFFFFFFF0;
    // rom_array[18159] = 32'hFFFFFFF1;
    // rom_array[18160] = 32'hFFFFFFF1;
    // rom_array[18161] = 32'hFFFFFFF0;
    // rom_array[18162] = 32'hFFFFFFF0;
    // rom_array[18163] = 32'hFFFFFFF1;
    // rom_array[18164] = 32'hFFFFFFF1;
    // rom_array[18165] = 32'hFFFFFFF0;
    // rom_array[18166] = 32'hFFFFFFF0;
    // rom_array[18167] = 32'hFFFFFFF1;
    // rom_array[18168] = 32'hFFFFFFF1;
    // rom_array[18169] = 32'hFFFFFFF0;
    // rom_array[18170] = 32'hFFFFFFF0;
    // rom_array[18171] = 32'hFFFFFFF1;
    // rom_array[18172] = 32'hFFFFFFF1;
    // rom_array[18173] = 32'hFFFFFFF0;
    // rom_array[18174] = 32'hFFFFFFF0;
    // rom_array[18175] = 32'hFFFFFFF0;
    // rom_array[18176] = 32'hFFFFFFF0;
    // rom_array[18177] = 32'hFFFFFFF0;
    // rom_array[18178] = 32'hFFFFFFF0;
    // rom_array[18179] = 32'hFFFFFFF1;
    // rom_array[18180] = 32'hFFFFFFF1;
    // rom_array[18181] = 32'hFFFFFFF0;
    // rom_array[18182] = 32'hFFFFFFF0;
    // rom_array[18183] = 32'hFFFFFFF0;
    // rom_array[18184] = 32'hFFFFFFF0;
    // rom_array[18185] = 32'hFFFFFFF1;
    // rom_array[18186] = 32'hFFFFFFF1;
    // rom_array[18187] = 32'hFFFFFFF1;
    // rom_array[18188] = 32'hFFFFFFF1;
    // rom_array[18189] = 32'hFFFFFFF0;
    // rom_array[18190] = 32'hFFFFFFF0;
    // rom_array[18191] = 32'hFFFFFFF0;
    // rom_array[18192] = 32'hFFFFFFF0;
    // rom_array[18193] = 32'hFFFFFFF1;
    // rom_array[18194] = 32'hFFFFFFF1;
    // rom_array[18195] = 32'hFFFFFFF1;
    // rom_array[18196] = 32'hFFFFFFF1;
    // rom_array[18197] = 32'hFFFFFFF0;
    // rom_array[18198] = 32'hFFFFFFF0;
    // rom_array[18199] = 32'hFFFFFFF0;
    // rom_array[18200] = 32'hFFFFFFF0;
    // rom_array[18201] = 32'hFFFFFFF1;
    // rom_array[18202] = 32'hFFFFFFF1;
    // rom_array[18203] = 32'hFFFFFFF1;
    // rom_array[18204] = 32'hFFFFFFF1;
    // rom_array[18205] = 32'hFFFFFFF0;
    // rom_array[18206] = 32'hFFFFFFF0;
    // rom_array[18207] = 32'hFFFFFFF0;
    // rom_array[18208] = 32'hFFFFFFF0;
    // rom_array[18209] = 32'hFFFFFFF1;
    // rom_array[18210] = 32'hFFFFFFF1;
    // rom_array[18211] = 32'hFFFFFFF1;
    // rom_array[18212] = 32'hFFFFFFF1;
    // rom_array[18213] = 32'hFFFFFFF0;
    // rom_array[18214] = 32'hFFFFFFF0;
    // rom_array[18215] = 32'hFFFFFFF0;
    // rom_array[18216] = 32'hFFFFFFF0;
    // rom_array[18217] = 32'hFFFFFFF1;
    // rom_array[18218] = 32'hFFFFFFF1;
    // rom_array[18219] = 32'hFFFFFFF1;
    // rom_array[18220] = 32'hFFFFFFF1;
    // rom_array[18221] = 32'hFFFFFFF0;
    // rom_array[18222] = 32'hFFFFFFF0;
    // rom_array[18223] = 32'hFFFFFFF0;
    // rom_array[18224] = 32'hFFFFFFF0;
    // rom_array[18225] = 32'hFFFFFFF1;
    // rom_array[18226] = 32'hFFFFFFF1;
    // rom_array[18227] = 32'hFFFFFFF1;
    // rom_array[18228] = 32'hFFFFFFF1;
    // rom_array[18229] = 32'hFFFFFFF0;
    // rom_array[18230] = 32'hFFFFFFF0;
    // rom_array[18231] = 32'hFFFFFFF0;
    // rom_array[18232] = 32'hFFFFFFF0;
    // rom_array[18233] = 32'hFFFFFFF1;
    // rom_array[18234] = 32'hFFFFFFF1;
    // rom_array[18235] = 32'hFFFFFFF1;
    // rom_array[18236] = 32'hFFFFFFF1;
    // rom_array[18237] = 32'hFFFFFFF1;
    // rom_array[18238] = 32'hFFFFFFF1;
    // rom_array[18239] = 32'hFFFFFFF1;
    // rom_array[18240] = 32'hFFFFFFF1;
    // rom_array[18241] = 32'hFFFFFFF1;
    // rom_array[18242] = 32'hFFFFFFF1;
    // rom_array[18243] = 32'hFFFFFFF1;
    // rom_array[18244] = 32'hFFFFFFF1;
    // rom_array[18245] = 32'hFFFFFFF1;
    // rom_array[18246] = 32'hFFFFFFF1;
    // rom_array[18247] = 32'hFFFFFFF1;
    // rom_array[18248] = 32'hFFFFFFF1;
    // rom_array[18249] = 32'hFFFFFFF1;
    // rom_array[18250] = 32'hFFFFFFF1;
    // rom_array[18251] = 32'hFFFFFFF1;
    // rom_array[18252] = 32'hFFFFFFF1;
    // rom_array[18253] = 32'hFFFFFFF1;
    // rom_array[18254] = 32'hFFFFFFF1;
    // rom_array[18255] = 32'hFFFFFFF1;
    // rom_array[18256] = 32'hFFFFFFF1;
    // rom_array[18257] = 32'hFFFFFFF1;
    // rom_array[18258] = 32'hFFFFFFF1;
    // rom_array[18259] = 32'hFFFFFFF1;
    // rom_array[18260] = 32'hFFFFFFF1;
    // rom_array[18261] = 32'hFFFFFFF1;
    // rom_array[18262] = 32'hFFFFFFF1;
    // rom_array[18263] = 32'hFFFFFFF1;
    // rom_array[18264] = 32'hFFFFFFF1;
    // rom_array[18265] = 32'hFFFFFFF1;
    // rom_array[18266] = 32'hFFFFFFF1;
    // rom_array[18267] = 32'hFFFFFFF1;
    // rom_array[18268] = 32'hFFFFFFF1;
    // rom_array[18269] = 32'hFFFFFFF0;
    // rom_array[18270] = 32'hFFFFFFF0;
    // rom_array[18271] = 32'hFFFFFFF0;
    // rom_array[18272] = 32'hFFFFFFF0;
    // rom_array[18273] = 32'hFFFFFFF1;
    // rom_array[18274] = 32'hFFFFFFF1;
    // rom_array[18275] = 32'hFFFFFFF1;
    // rom_array[18276] = 32'hFFFFFFF1;
    // rom_array[18277] = 32'hFFFFFFF0;
    // rom_array[18278] = 32'hFFFFFFF0;
    // rom_array[18279] = 32'hFFFFFFF0;
    // rom_array[18280] = 32'hFFFFFFF0;
    // rom_array[18281] = 32'hFFFFFFF1;
    // rom_array[18282] = 32'hFFFFFFF1;
    // rom_array[18283] = 32'hFFFFFFF1;
    // rom_array[18284] = 32'hFFFFFFF1;
    // rom_array[18285] = 32'hFFFFFFF0;
    // rom_array[18286] = 32'hFFFFFFF0;
    // rom_array[18287] = 32'hFFFFFFF0;
    // rom_array[18288] = 32'hFFFFFFF0;
    // rom_array[18289] = 32'hFFFFFFF1;
    // rom_array[18290] = 32'hFFFFFFF1;
    // rom_array[18291] = 32'hFFFFFFF1;
    // rom_array[18292] = 32'hFFFFFFF1;
    // rom_array[18293] = 32'hFFFFFFF0;
    // rom_array[18294] = 32'hFFFFFFF0;
    // rom_array[18295] = 32'hFFFFFFF0;
    // rom_array[18296] = 32'hFFFFFFF0;
    // rom_array[18297] = 32'hFFFFFFF1;
    // rom_array[18298] = 32'hFFFFFFF1;
    // rom_array[18299] = 32'hFFFFFFF1;
    // rom_array[18300] = 32'hFFFFFFF1;
    // rom_array[18301] = 32'hFFFFFFF0;
    // rom_array[18302] = 32'hFFFFFFF0;
    // rom_array[18303] = 32'hFFFFFFF0;
    // rom_array[18304] = 32'hFFFFFFF0;
    // rom_array[18305] = 32'hFFFFFFF1;
    // rom_array[18306] = 32'hFFFFFFF1;
    // rom_array[18307] = 32'hFFFFFFF1;
    // rom_array[18308] = 32'hFFFFFFF1;
    // rom_array[18309] = 32'hFFFFFFF0;
    // rom_array[18310] = 32'hFFFFFFF0;
    // rom_array[18311] = 32'hFFFFFFF0;
    // rom_array[18312] = 32'hFFFFFFF0;
    // rom_array[18313] = 32'hFFFFFFF1;
    // rom_array[18314] = 32'hFFFFFFF1;
    // rom_array[18315] = 32'hFFFFFFF1;
    // rom_array[18316] = 32'hFFFFFFF1;
    // rom_array[18317] = 32'hFFFFFFF1;
    // rom_array[18318] = 32'hFFFFFFF1;
    // rom_array[18319] = 32'hFFFFFFF1;
    // rom_array[18320] = 32'hFFFFFFF1;
    // rom_array[18321] = 32'hFFFFFFF1;
    // rom_array[18322] = 32'hFFFFFFF1;
    // rom_array[18323] = 32'hFFFFFFF1;
    // rom_array[18324] = 32'hFFFFFFF1;
    // rom_array[18325] = 32'hFFFFFFF1;
    // rom_array[18326] = 32'hFFFFFFF1;
    // rom_array[18327] = 32'hFFFFFFF1;
    // rom_array[18328] = 32'hFFFFFFF1;
    // rom_array[18329] = 32'hFFFFFFF1;
    // rom_array[18330] = 32'hFFFFFFF1;
    // rom_array[18331] = 32'hFFFFFFF1;
    // rom_array[18332] = 32'hFFFFFFF1;
    // rom_array[18333] = 32'hFFFFFFF1;
    // rom_array[18334] = 32'hFFFFFFF1;
    // rom_array[18335] = 32'hFFFFFFF1;
    // rom_array[18336] = 32'hFFFFFFF1;
    // rom_array[18337] = 32'hFFFFFFF1;
    // rom_array[18338] = 32'hFFFFFFF1;
    // rom_array[18339] = 32'hFFFFFFF1;
    // rom_array[18340] = 32'hFFFFFFF1;
    // rom_array[18341] = 32'hFFFFFFF1;
    // rom_array[18342] = 32'hFFFFFFF1;
    // rom_array[18343] = 32'hFFFFFFF1;
    // rom_array[18344] = 32'hFFFFFFF1;
    // rom_array[18345] = 32'hFFFFFFF1;
    // rom_array[18346] = 32'hFFFFFFF1;
    // rom_array[18347] = 32'hFFFFFFF1;
    // rom_array[18348] = 32'hFFFFFFF1;
    // rom_array[18349] = 32'hFFFFFFF0;
    // rom_array[18350] = 32'hFFFFFFF0;
    // rom_array[18351] = 32'hFFFFFFF0;
    // rom_array[18352] = 32'hFFFFFFF0;
    // rom_array[18353] = 32'hFFFFFFF1;
    // rom_array[18354] = 32'hFFFFFFF1;
    // rom_array[18355] = 32'hFFFFFFF1;
    // rom_array[18356] = 32'hFFFFFFF1;
    // rom_array[18357] = 32'hFFFFFFF0;
    // rom_array[18358] = 32'hFFFFFFF0;
    // rom_array[18359] = 32'hFFFFFFF0;
    // rom_array[18360] = 32'hFFFFFFF0;
    // rom_array[18361] = 32'hFFFFFFF1;
    // rom_array[18362] = 32'hFFFFFFF1;
    // rom_array[18363] = 32'hFFFFFFF1;
    // rom_array[18364] = 32'hFFFFFFF1;
    // rom_array[18365] = 32'hFFFFFFF0;
    // rom_array[18366] = 32'hFFFFFFF0;
    // rom_array[18367] = 32'hFFFFFFF0;
    // rom_array[18368] = 32'hFFFFFFF0;
    // rom_array[18369] = 32'hFFFFFFF1;
    // rom_array[18370] = 32'hFFFFFFF1;
    // rom_array[18371] = 32'hFFFFFFF1;
    // rom_array[18372] = 32'hFFFFFFF1;
    // rom_array[18373] = 32'hFFFFFFF0;
    // rom_array[18374] = 32'hFFFFFFF0;
    // rom_array[18375] = 32'hFFFFFFF0;
    // rom_array[18376] = 32'hFFFFFFF0;
    // rom_array[18377] = 32'hFFFFFFF1;
    // rom_array[18378] = 32'hFFFFFFF1;
    // rom_array[18379] = 32'hFFFFFFF1;
    // rom_array[18380] = 32'hFFFFFFF1;
    // rom_array[18381] = 32'hFFFFFFF0;
    // rom_array[18382] = 32'hFFFFFFF0;
    // rom_array[18383] = 32'hFFFFFFF0;
    // rom_array[18384] = 32'hFFFFFFF0;
    // rom_array[18385] = 32'hFFFFFFF1;
    // rom_array[18386] = 32'hFFFFFFF1;
    // rom_array[18387] = 32'hFFFFFFF1;
    // rom_array[18388] = 32'hFFFFFFF1;
    // rom_array[18389] = 32'hFFFFFFF0;
    // rom_array[18390] = 32'hFFFFFFF0;
    // rom_array[18391] = 32'hFFFFFFF0;
    // rom_array[18392] = 32'hFFFFFFF0;
    // rom_array[18393] = 32'hFFFFFFF1;
    // rom_array[18394] = 32'hFFFFFFF1;
    // rom_array[18395] = 32'hFFFFFFF1;
    // rom_array[18396] = 32'hFFFFFFF1;
    // rom_array[18397] = 32'hFFFFFFF0;
    // rom_array[18398] = 32'hFFFFFFF0;
    // rom_array[18399] = 32'hFFFFFFF0;
    // rom_array[18400] = 32'hFFFFFFF0;
    // rom_array[18401] = 32'hFFFFFFF1;
    // rom_array[18402] = 32'hFFFFFFF1;
    // rom_array[18403] = 32'hFFFFFFF1;
    // rom_array[18404] = 32'hFFFFFFF1;
    // rom_array[18405] = 32'hFFFFFFF0;
    // rom_array[18406] = 32'hFFFFFFF0;
    // rom_array[18407] = 32'hFFFFFFF0;
    // rom_array[18408] = 32'hFFFFFFF0;
    // rom_array[18409] = 32'hFFFFFFF1;
    // rom_array[18410] = 32'hFFFFFFF1;
    // rom_array[18411] = 32'hFFFFFFF1;
    // rom_array[18412] = 32'hFFFFFFF1;
    // rom_array[18413] = 32'hFFFFFFF1;
    // rom_array[18414] = 32'hFFFFFFF1;
    // rom_array[18415] = 32'hFFFFFFF1;
    // rom_array[18416] = 32'hFFFFFFF1;
    // rom_array[18417] = 32'hFFFFFFF1;
    // rom_array[18418] = 32'hFFFFFFF1;
    // rom_array[18419] = 32'hFFFFFFF1;
    // rom_array[18420] = 32'hFFFFFFF1;
    // rom_array[18421] = 32'hFFFFFFF1;
    // rom_array[18422] = 32'hFFFFFFF1;
    // rom_array[18423] = 32'hFFFFFFF1;
    // rom_array[18424] = 32'hFFFFFFF1;
    // rom_array[18425] = 32'hFFFFFFF1;
    // rom_array[18426] = 32'hFFFFFFF1;
    // rom_array[18427] = 32'hFFFFFFF1;
    // rom_array[18428] = 32'hFFFFFFF1;
    // rom_array[18429] = 32'hFFFFFFF1;
    // rom_array[18430] = 32'hFFFFFFF1;
    // rom_array[18431] = 32'hFFFFFFF1;
    // rom_array[18432] = 32'hFFFFFFF1;
    // rom_array[18433] = 32'hFFFFFFF1;
    // rom_array[18434] = 32'hFFFFFFF1;
    // rom_array[18435] = 32'hFFFFFFF1;
    // rom_array[18436] = 32'hFFFFFFF1;
    // rom_array[18437] = 32'hFFFFFFF1;
    // rom_array[18438] = 32'hFFFFFFF1;
    // rom_array[18439] = 32'hFFFFFFF1;
    // rom_array[18440] = 32'hFFFFFFF1;
    // rom_array[18441] = 32'hFFFFFFF1;
    // rom_array[18442] = 32'hFFFFFFF1;
    // rom_array[18443] = 32'hFFFFFFF1;
    // rom_array[18444] = 32'hFFFFFFF1;
    // rom_array[18445] = 32'hFFFFFFF1;
    // rom_array[18446] = 32'hFFFFFFF1;
    // rom_array[18447] = 32'hFFFFFFF1;
    // rom_array[18448] = 32'hFFFFFFF1;
    // rom_array[18449] = 32'hFFFFFFF1;
    // rom_array[18450] = 32'hFFFFFFF1;
    // rom_array[18451] = 32'hFFFFFFF1;
    // rom_array[18452] = 32'hFFFFFFF1;
    // rom_array[18453] = 32'hFFFFFFF1;
    // rom_array[18454] = 32'hFFFFFFF1;
    // rom_array[18455] = 32'hFFFFFFF1;
    // rom_array[18456] = 32'hFFFFFFF1;
    // rom_array[18457] = 32'hFFFFFFF1;
    // rom_array[18458] = 32'hFFFFFFF1;
    // rom_array[18459] = 32'hFFFFFFF1;
    // rom_array[18460] = 32'hFFFFFFF1;
    // rom_array[18461] = 32'hFFFFFFF1;
    // rom_array[18462] = 32'hFFFFFFF1;
    // rom_array[18463] = 32'hFFFFFFF1;
    // rom_array[18464] = 32'hFFFFFFF1;
    // rom_array[18465] = 32'hFFFFFFF1;
    // rom_array[18466] = 32'hFFFFFFF1;
    // rom_array[18467] = 32'hFFFFFFF1;
    // rom_array[18468] = 32'hFFFFFFF1;
    // rom_array[18469] = 32'hFFFFFFF1;
    // rom_array[18470] = 32'hFFFFFFF1;
    // rom_array[18471] = 32'hFFFFFFF1;
    // rom_array[18472] = 32'hFFFFFFF1;
    // rom_array[18473] = 32'hFFFFFFF1;
    // rom_array[18474] = 32'hFFFFFFF1;
    // rom_array[18475] = 32'hFFFFFFF1;
    // rom_array[18476] = 32'hFFFFFFF1;
    // rom_array[18477] = 32'hFFFFFFF1;
    // rom_array[18478] = 32'hFFFFFFF1;
    // rom_array[18479] = 32'hFFFFFFF1;
    // rom_array[18480] = 32'hFFFFFFF1;
    // rom_array[18481] = 32'hFFFFFFF1;
    // rom_array[18482] = 32'hFFFFFFF1;
    // rom_array[18483] = 32'hFFFFFFF1;
    // rom_array[18484] = 32'hFFFFFFF1;
    // rom_array[18485] = 32'hFFFFFFF1;
    // rom_array[18486] = 32'hFFFFFFF1;
    // rom_array[18487] = 32'hFFFFFFF1;
    // rom_array[18488] = 32'hFFFFFFF1;
    // rom_array[18489] = 32'hFFFFFFF1;
    // rom_array[18490] = 32'hFFFFFFF1;
    // rom_array[18491] = 32'hFFFFFFF1;
    // rom_array[18492] = 32'hFFFFFFF1;
    // rom_array[18493] = 32'hFFFFFFF1;
    // rom_array[18494] = 32'hFFFFFFF1;
    // rom_array[18495] = 32'hFFFFFFF1;
    // rom_array[18496] = 32'hFFFFFFF1;
    // rom_array[18497] = 32'hFFFFFFF1;
    // rom_array[18498] = 32'hFFFFFFF1;
    // rom_array[18499] = 32'hFFFFFFF1;
    // rom_array[18500] = 32'hFFFFFFF1;
    // rom_array[18501] = 32'hFFFFFFF1;
    // rom_array[18502] = 32'hFFFFFFF1;
    // rom_array[18503] = 32'hFFFFFFF1;
    // rom_array[18504] = 32'hFFFFFFF1;
    // rom_array[18505] = 32'hFFFFFFF1;
    // rom_array[18506] = 32'hFFFFFFF1;
    // rom_array[18507] = 32'hFFFFFFF1;
    // rom_array[18508] = 32'hFFFFFFF1;
    // rom_array[18509] = 32'hFFFFFFF1;
    // rom_array[18510] = 32'hFFFFFFF1;
    // rom_array[18511] = 32'hFFFFFFF1;
    // rom_array[18512] = 32'hFFFFFFF1;
    // rom_array[18513] = 32'hFFFFFFF1;
    // rom_array[18514] = 32'hFFFFFFF1;
    // rom_array[18515] = 32'hFFFFFFF1;
    // rom_array[18516] = 32'hFFFFFFF1;
    // rom_array[18517] = 32'hFFFFFFF1;
    // rom_array[18518] = 32'hFFFFFFF1;
    // rom_array[18519] = 32'hFFFFFFF1;
    // rom_array[18520] = 32'hFFFFFFF1;
    // rom_array[18521] = 32'hFFFFFFF1;
    // rom_array[18522] = 32'hFFFFFFF1;
    // rom_array[18523] = 32'hFFFFFFF1;
    // rom_array[18524] = 32'hFFFFFFF1;
    // rom_array[18525] = 32'hFFFFFFF1;
    // rom_array[18526] = 32'hFFFFFFF1;
    // rom_array[18527] = 32'hFFFFFFF1;
    // rom_array[18528] = 32'hFFFFFFF1;
    // rom_array[18529] = 32'hFFFFFFF1;
    // rom_array[18530] = 32'hFFFFFFF1;
    // rom_array[18531] = 32'hFFFFFFF1;
    // rom_array[18532] = 32'hFFFFFFF1;
    // rom_array[18533] = 32'hFFFFFFF1;
    // rom_array[18534] = 32'hFFFFFFF1;
    // rom_array[18535] = 32'hFFFFFFF1;
    // rom_array[18536] = 32'hFFFFFFF1;
    // rom_array[18537] = 32'hFFFFFFF1;
    // rom_array[18538] = 32'hFFFFFFF1;
    // rom_array[18539] = 32'hFFFFFFF1;
    // rom_array[18540] = 32'hFFFFFFF1;
    // rom_array[18541] = 32'hFFFFFFF1;
    // rom_array[18542] = 32'hFFFFFFF1;
    // rom_array[18543] = 32'hFFFFFFF1;
    // rom_array[18544] = 32'hFFFFFFF1;
    // rom_array[18545] = 32'hFFFFFFF1;
    // rom_array[18546] = 32'hFFFFFFF1;
    // rom_array[18547] = 32'hFFFFFFF1;
    // rom_array[18548] = 32'hFFFFFFF1;
    // rom_array[18549] = 32'hFFFFFFF1;
    // rom_array[18550] = 32'hFFFFFFF1;
    // rom_array[18551] = 32'hFFFFFFF1;
    // rom_array[18552] = 32'hFFFFFFF1;
    // rom_array[18553] = 32'hFFFFFFF1;
    // rom_array[18554] = 32'hFFFFFFF1;
    // rom_array[18555] = 32'hFFFFFFF1;
    // rom_array[18556] = 32'hFFFFFFF1;
    // rom_array[18557] = 32'hFFFFFFF1;
    // rom_array[18558] = 32'hFFFFFFF1;
    // rom_array[18559] = 32'hFFFFFFF1;
    // rom_array[18560] = 32'hFFFFFFF1;
    // rom_array[18561] = 32'hFFFFFFF1;
    // rom_array[18562] = 32'hFFFFFFF1;
    // rom_array[18563] = 32'hFFFFFFF1;
    // rom_array[18564] = 32'hFFFFFFF1;
    // rom_array[18565] = 32'hFFFFFFF1;
    // rom_array[18566] = 32'hFFFFFFF1;
    // rom_array[18567] = 32'hFFFFFFF1;
    // rom_array[18568] = 32'hFFFFFFF1;
    // rom_array[18569] = 32'hFFFFFFF1;
    // rom_array[18570] = 32'hFFFFFFF1;
    // rom_array[18571] = 32'hFFFFFFF1;
    // rom_array[18572] = 32'hFFFFFFF1;
    // rom_array[18573] = 32'hFFFFFFF1;
    // rom_array[18574] = 32'hFFFFFFF1;
    // rom_array[18575] = 32'hFFFFFFF1;
    // rom_array[18576] = 32'hFFFFFFF1;
    // rom_array[18577] = 32'hFFFFFFF1;
    // rom_array[18578] = 32'hFFFFFFF1;
    // rom_array[18579] = 32'hFFFFFFF1;
    // rom_array[18580] = 32'hFFFFFFF1;
    // rom_array[18581] = 32'hFFFFFFF1;
    // rom_array[18582] = 32'hFFFFFFF1;
    // rom_array[18583] = 32'hFFFFFFF1;
    // rom_array[18584] = 32'hFFFFFFF1;
    // rom_array[18585] = 32'hFFFFFFF1;
    // rom_array[18586] = 32'hFFFFFFF1;
    // rom_array[18587] = 32'hFFFFFFF1;
    // rom_array[18588] = 32'hFFFFFFF1;
    // rom_array[18589] = 32'hFFFFFFF1;
    // rom_array[18590] = 32'hFFFFFFF1;
    // rom_array[18591] = 32'hFFFFFFF1;
    // rom_array[18592] = 32'hFFFFFFF1;
    // rom_array[18593] = 32'hFFFFFFF1;
    // rom_array[18594] = 32'hFFFFFFF1;
    // rom_array[18595] = 32'hFFFFFFF1;
    // rom_array[18596] = 32'hFFFFFFF1;
    // rom_array[18597] = 32'hFFFFFFF1;
    // rom_array[18598] = 32'hFFFFFFF1;
    // rom_array[18599] = 32'hFFFFFFF1;
    // rom_array[18600] = 32'hFFFFFFF1;
    // rom_array[18601] = 32'hFFFFFFF1;
    // rom_array[18602] = 32'hFFFFFFF1;
    // rom_array[18603] = 32'hFFFFFFF1;
    // rom_array[18604] = 32'hFFFFFFF1;
    // rom_array[18605] = 32'hFFFFFFF1;
    // rom_array[18606] = 32'hFFFFFFF1;
    // rom_array[18607] = 32'hFFFFFFF1;
    // rom_array[18608] = 32'hFFFFFFF1;
    // rom_array[18609] = 32'hFFFFFFF1;
    // rom_array[18610] = 32'hFFFFFFF1;
    // rom_array[18611] = 32'hFFFFFFF1;
    // rom_array[18612] = 32'hFFFFFFF1;
    // rom_array[18613] = 32'hFFFFFFF1;
    // rom_array[18614] = 32'hFFFFFFF1;
    // rom_array[18615] = 32'hFFFFFFF1;
    // rom_array[18616] = 32'hFFFFFFF1;
    // rom_array[18617] = 32'hFFFFFFF1;
    // rom_array[18618] = 32'hFFFFFFF1;
    // rom_array[18619] = 32'hFFFFFFF1;
    // rom_array[18620] = 32'hFFFFFFF1;
    // rom_array[18621] = 32'hFFFFFFF1;
    // rom_array[18622] = 32'hFFFFFFF1;
    // rom_array[18623] = 32'hFFFFFFF1;
    // rom_array[18624] = 32'hFFFFFFF1;
    // rom_array[18625] = 32'hFFFFFFF1;
    // rom_array[18626] = 32'hFFFFFFF1;
    // rom_array[18627] = 32'hFFFFFFF1;
    // rom_array[18628] = 32'hFFFFFFF1;
    // rom_array[18629] = 32'hFFFFFFF1;
    // rom_array[18630] = 32'hFFFFFFF1;
    // rom_array[18631] = 32'hFFFFFFF1;
    // rom_array[18632] = 32'hFFFFFFF1;
    // rom_array[18633] = 32'hFFFFFFF1;
    // rom_array[18634] = 32'hFFFFFFF1;
    // rom_array[18635] = 32'hFFFFFFF1;
    // rom_array[18636] = 32'hFFFFFFF1;
    // rom_array[18637] = 32'hFFFFFFF1;
    // rom_array[18638] = 32'hFFFFFFF1;
    // rom_array[18639] = 32'hFFFFFFF1;
    // rom_array[18640] = 32'hFFFFFFF1;
    // rom_array[18641] = 32'hFFFFFFF1;
    // rom_array[18642] = 32'hFFFFFFF1;
    // rom_array[18643] = 32'hFFFFFFF1;
    // rom_array[18644] = 32'hFFFFFFF1;
    // rom_array[18645] = 32'hFFFFFFF1;
    // rom_array[18646] = 32'hFFFFFFF1;
    // rom_array[18647] = 32'hFFFFFFF1;
    // rom_array[18648] = 32'hFFFFFFF1;
    // rom_array[18649] = 32'hFFFFFFF1;
    // rom_array[18650] = 32'hFFFFFFF1;
    // rom_array[18651] = 32'hFFFFFFF1;
    // rom_array[18652] = 32'hFFFFFFF1;
    // rom_array[18653] = 32'hFFFFFFF1;
    // rom_array[18654] = 32'hFFFFFFF1;
    // rom_array[18655] = 32'hFFFFFFF1;
    // rom_array[18656] = 32'hFFFFFFF1;
    // rom_array[18657] = 32'hFFFFFFF1;
    // rom_array[18658] = 32'hFFFFFFF1;
    // rom_array[18659] = 32'hFFFFFFF1;
    // rom_array[18660] = 32'hFFFFFFF1;
    // rom_array[18661] = 32'hFFFFFFF1;
    // rom_array[18662] = 32'hFFFFFFF1;
    // rom_array[18663] = 32'hFFFFFFF1;
    // rom_array[18664] = 32'hFFFFFFF1;
    // rom_array[18665] = 32'hFFFFFFF1;
    // rom_array[18666] = 32'hFFFFFFF1;
    // rom_array[18667] = 32'hFFFFFFF1;
    // rom_array[18668] = 32'hFFFFFFF1;
    // rom_array[18669] = 32'hFFFFFFF1;
    // rom_array[18670] = 32'hFFFFFFF1;
    // rom_array[18671] = 32'hFFFFFFF1;
    // rom_array[18672] = 32'hFFFFFFF1;
    // rom_array[18673] = 32'hFFFFFFF1;
    // rom_array[18674] = 32'hFFFFFFF1;
    // rom_array[18675] = 32'hFFFFFFF1;
    // rom_array[18676] = 32'hFFFFFFF1;
    // rom_array[18677] = 32'hFFFFFFF1;
    // rom_array[18678] = 32'hFFFFFFF1;
    // rom_array[18679] = 32'hFFFFFFF1;
    // rom_array[18680] = 32'hFFFFFFF1;
    // rom_array[18681] = 32'hFFFFFFF1;
    // rom_array[18682] = 32'hFFFFFFF1;
    // rom_array[18683] = 32'hFFFFFFF1;
    // rom_array[18684] = 32'hFFFFFFF1;
    // rom_array[18685] = 32'hFFFFFFF1;
    // rom_array[18686] = 32'hFFFFFFF1;
    // rom_array[18687] = 32'hFFFFFFF1;
    // rom_array[18688] = 32'hFFFFFFF1;
    // rom_array[18689] = 32'hFFFFFFF1;
    // rom_array[18690] = 32'hFFFFFFF1;
    // rom_array[18691] = 32'hFFFFFFF1;
    // rom_array[18692] = 32'hFFFFFFF1;
    // rom_array[18693] = 32'hFFFFFFF1;
    // rom_array[18694] = 32'hFFFFFFF1;
    // rom_array[18695] = 32'hFFFFFFF1;
    // rom_array[18696] = 32'hFFFFFFF1;
    // rom_array[18697] = 32'hFFFFFFF1;
    // rom_array[18698] = 32'hFFFFFFF1;
    // rom_array[18699] = 32'hFFFFFFF1;
    // rom_array[18700] = 32'hFFFFFFF1;
    // rom_array[18701] = 32'hFFFFFFF1;
    // rom_array[18702] = 32'hFFFFFFF1;
    // rom_array[18703] = 32'hFFFFFFF1;
    // rom_array[18704] = 32'hFFFFFFF1;
    // rom_array[18705] = 32'hFFFFFFF1;
    // rom_array[18706] = 32'hFFFFFFF1;
    // rom_array[18707] = 32'hFFFFFFF1;
    // rom_array[18708] = 32'hFFFFFFF1;
    // rom_array[18709] = 32'hFFFFFFF1;
    // rom_array[18710] = 32'hFFFFFFF1;
    // rom_array[18711] = 32'hFFFFFFF1;
    // rom_array[18712] = 32'hFFFFFFF1;
    // rom_array[18713] = 32'hFFFFFFF1;
    // rom_array[18714] = 32'hFFFFFFF1;
    // rom_array[18715] = 32'hFFFFFFF1;
    // rom_array[18716] = 32'hFFFFFFF1;
    // rom_array[18717] = 32'hFFFFFFF1;
    // rom_array[18718] = 32'hFFFFFFF1;
    // rom_array[18719] = 32'hFFFFFFF1;
    // rom_array[18720] = 32'hFFFFFFF1;
    // rom_array[18721] = 32'hFFFFFFF1;
    // rom_array[18722] = 32'hFFFFFFF1;
    // rom_array[18723] = 32'hFFFFFFF1;
    // rom_array[18724] = 32'hFFFFFFF1;
    // rom_array[18725] = 32'hFFFFFFF1;
    // rom_array[18726] = 32'hFFFFFFF1;
    // rom_array[18727] = 32'hFFFFFFF1;
    // rom_array[18728] = 32'hFFFFFFF1;
    // rom_array[18729] = 32'hFFFFFFF1;
    // rom_array[18730] = 32'hFFFFFFF1;
    // rom_array[18731] = 32'hFFFFFFF1;
    // rom_array[18732] = 32'hFFFFFFF1;
    // rom_array[18733] = 32'hFFFFFFF1;
    // rom_array[18734] = 32'hFFFFFFF1;
    // rom_array[18735] = 32'hFFFFFFF1;
    // rom_array[18736] = 32'hFFFFFFF1;
    // rom_array[18737] = 32'hFFFFFFF1;
    // rom_array[18738] = 32'hFFFFFFF1;
    // rom_array[18739] = 32'hFFFFFFF1;
    // rom_array[18740] = 32'hFFFFFFF1;
    // rom_array[18741] = 32'hFFFFFFF1;
    // rom_array[18742] = 32'hFFFFFFF1;
    // rom_array[18743] = 32'hFFFFFFF1;
    // rom_array[18744] = 32'hFFFFFFF1;
    // rom_array[18745] = 32'hFFFFFFF1;
    // rom_array[18746] = 32'hFFFFFFF1;
    // rom_array[18747] = 32'hFFFFFFF1;
    // rom_array[18748] = 32'hFFFFFFF1;
    // rom_array[18749] = 32'hFFFFFFF1;
    // rom_array[18750] = 32'hFFFFFFF1;
    // rom_array[18751] = 32'hFFFFFFF1;
    // rom_array[18752] = 32'hFFFFFFF1;
    // rom_array[18753] = 32'hFFFFFFF1;
    // rom_array[18754] = 32'hFFFFFFF1;
    // rom_array[18755] = 32'hFFFFFFF1;
    // rom_array[18756] = 32'hFFFFFFF1;
    // rom_array[18757] = 32'hFFFFFFF1;
    // rom_array[18758] = 32'hFFFFFFF1;
    // rom_array[18759] = 32'hFFFFFFF1;
    // rom_array[18760] = 32'hFFFFFFF1;
    // rom_array[18761] = 32'hFFFFFFF1;
    // rom_array[18762] = 32'hFFFFFFF1;
    // rom_array[18763] = 32'hFFFFFFF1;
    // rom_array[18764] = 32'hFFFFFFF1;
    // rom_array[18765] = 32'hFFFFFFF1;
    // rom_array[18766] = 32'hFFFFFFF1;
    // rom_array[18767] = 32'hFFFFFFF1;
    // rom_array[18768] = 32'hFFFFFFF1;
    // rom_array[18769] = 32'hFFFFFFF1;
    // rom_array[18770] = 32'hFFFFFFF1;
    // rom_array[18771] = 32'hFFFFFFF1;
    // rom_array[18772] = 32'hFFFFFFF1;
    // rom_array[18773] = 32'hFFFFFFF1;
    // rom_array[18774] = 32'hFFFFFFF1;
    // rom_array[18775] = 32'hFFFFFFF1;
    // rom_array[18776] = 32'hFFFFFFF1;
    // rom_array[18777] = 32'hFFFFFFF0;
    // rom_array[18778] = 32'hFFFFFFF0;
    // rom_array[18779] = 32'hFFFFFFF0;
    // rom_array[18780] = 32'hFFFFFFF0;
    // rom_array[18781] = 32'hFFFFFFF0;
    // rom_array[18782] = 32'hFFFFFFF0;
    // rom_array[18783] = 32'hFFFFFFF1;
    // rom_array[18784] = 32'hFFFFFFF1;
    // rom_array[18785] = 32'hFFFFFFF0;
    // rom_array[18786] = 32'hFFFFFFF0;
    // rom_array[18787] = 32'hFFFFFFF0;
    // rom_array[18788] = 32'hFFFFFFF0;
    // rom_array[18789] = 32'hFFFFFFF0;
    // rom_array[18790] = 32'hFFFFFFF0;
    // rom_array[18791] = 32'hFFFFFFF1;
    // rom_array[18792] = 32'hFFFFFFF1;
    // rom_array[18793] = 32'hFFFFFFF0;
    // rom_array[18794] = 32'hFFFFFFF0;
    // rom_array[18795] = 32'hFFFFFFF0;
    // rom_array[18796] = 32'hFFFFFFF0;
    // rom_array[18797] = 32'hFFFFFFF1;
    // rom_array[18798] = 32'hFFFFFFF1;
    // rom_array[18799] = 32'hFFFFFFF1;
    // rom_array[18800] = 32'hFFFFFFF1;
    // rom_array[18801] = 32'hFFFFFFF0;
    // rom_array[18802] = 32'hFFFFFFF0;
    // rom_array[18803] = 32'hFFFFFFF0;
    // rom_array[18804] = 32'hFFFFFFF0;
    // rom_array[18805] = 32'hFFFFFFF1;
    // rom_array[18806] = 32'hFFFFFFF1;
    // rom_array[18807] = 32'hFFFFFFF1;
    // rom_array[18808] = 32'hFFFFFFF1;
    // rom_array[18809] = 32'hFFFFFFF0;
    // rom_array[18810] = 32'hFFFFFFF0;
    // rom_array[18811] = 32'hFFFFFFF1;
    // rom_array[18812] = 32'hFFFFFFF1;
    // rom_array[18813] = 32'hFFFFFFF0;
    // rom_array[18814] = 32'hFFFFFFF0;
    // rom_array[18815] = 32'hFFFFFFF1;
    // rom_array[18816] = 32'hFFFFFFF1;
    // rom_array[18817] = 32'hFFFFFFF0;
    // rom_array[18818] = 32'hFFFFFFF0;
    // rom_array[18819] = 32'hFFFFFFF1;
    // rom_array[18820] = 32'hFFFFFFF1;
    // rom_array[18821] = 32'hFFFFFFF0;
    // rom_array[18822] = 32'hFFFFFFF0;
    // rom_array[18823] = 32'hFFFFFFF1;
    // rom_array[18824] = 32'hFFFFFFF1;
    // rom_array[18825] = 32'hFFFFFFF0;
    // rom_array[18826] = 32'hFFFFFFF0;
    // rom_array[18827] = 32'hFFFFFFF0;
    // rom_array[18828] = 32'hFFFFFFF0;
    // rom_array[18829] = 32'hFFFFFFF1;
    // rom_array[18830] = 32'hFFFFFFF1;
    // rom_array[18831] = 32'hFFFFFFF1;
    // rom_array[18832] = 32'hFFFFFFF1;
    // rom_array[18833] = 32'hFFFFFFF0;
    // rom_array[18834] = 32'hFFFFFFF0;
    // rom_array[18835] = 32'hFFFFFFF0;
    // rom_array[18836] = 32'hFFFFFFF0;
    // rom_array[18837] = 32'hFFFFFFF1;
    // rom_array[18838] = 32'hFFFFFFF1;
    // rom_array[18839] = 32'hFFFFFFF1;
    // rom_array[18840] = 32'hFFFFFFF1;
    // rom_array[18841] = 32'hFFFFFFF0;
    // rom_array[18842] = 32'hFFFFFFF0;
    // rom_array[18843] = 32'hFFFFFFF0;
    // rom_array[18844] = 32'hFFFFFFF0;
    // rom_array[18845] = 32'hFFFFFFF1;
    // rom_array[18846] = 32'hFFFFFFF1;
    // rom_array[18847] = 32'hFFFFFFF1;
    // rom_array[18848] = 32'hFFFFFFF1;
    // rom_array[18849] = 32'hFFFFFFF0;
    // rom_array[18850] = 32'hFFFFFFF0;
    // rom_array[18851] = 32'hFFFFFFF0;
    // rom_array[18852] = 32'hFFFFFFF0;
    // rom_array[18853] = 32'hFFFFFFF1;
    // rom_array[18854] = 32'hFFFFFFF1;
    // rom_array[18855] = 32'hFFFFFFF1;
    // rom_array[18856] = 32'hFFFFFFF1;
    // rom_array[18857] = 32'hFFFFFFF0;
    // rom_array[18858] = 32'hFFFFFFF0;
    // rom_array[18859] = 32'hFFFFFFF1;
    // rom_array[18860] = 32'hFFFFFFF1;
    // rom_array[18861] = 32'hFFFFFFF0;
    // rom_array[18862] = 32'hFFFFFFF0;
    // rom_array[18863] = 32'hFFFFFFF1;
    // rom_array[18864] = 32'hFFFFFFF1;
    // rom_array[18865] = 32'hFFFFFFF0;
    // rom_array[18866] = 32'hFFFFFFF0;
    // rom_array[18867] = 32'hFFFFFFF1;
    // rom_array[18868] = 32'hFFFFFFF1;
    // rom_array[18869] = 32'hFFFFFFF0;
    // rom_array[18870] = 32'hFFFFFFF0;
    // rom_array[18871] = 32'hFFFFFFF1;
    // rom_array[18872] = 32'hFFFFFFF1;
    // rom_array[18873] = 32'hFFFFFFF0;
    // rom_array[18874] = 32'hFFFFFFF0;
    // rom_array[18875] = 32'hFFFFFFF1;
    // rom_array[18876] = 32'hFFFFFFF1;
    // rom_array[18877] = 32'hFFFFFFF0;
    // rom_array[18878] = 32'hFFFFFFF0;
    // rom_array[18879] = 32'hFFFFFFF1;
    // rom_array[18880] = 32'hFFFFFFF1;
    // rom_array[18881] = 32'hFFFFFFF0;
    // rom_array[18882] = 32'hFFFFFFF0;
    // rom_array[18883] = 32'hFFFFFFF1;
    // rom_array[18884] = 32'hFFFFFFF1;
    // rom_array[18885] = 32'hFFFFFFF0;
    // rom_array[18886] = 32'hFFFFFFF0;
    // rom_array[18887] = 32'hFFFFFFF1;
    // rom_array[18888] = 32'hFFFFFFF1;
    // rom_array[18889] = 32'hFFFFFFF0;
    // rom_array[18890] = 32'hFFFFFFF0;
    // rom_array[18891] = 32'hFFFFFFF1;
    // rom_array[18892] = 32'hFFFFFFF1;
    // rom_array[18893] = 32'hFFFFFFF0;
    // rom_array[18894] = 32'hFFFFFFF0;
    // rom_array[18895] = 32'hFFFFFFF0;
    // rom_array[18896] = 32'hFFFFFFF0;
    // rom_array[18897] = 32'hFFFFFFF0;
    // rom_array[18898] = 32'hFFFFFFF0;
    // rom_array[18899] = 32'hFFFFFFF1;
    // rom_array[18900] = 32'hFFFFFFF1;
    // rom_array[18901] = 32'hFFFFFFF0;
    // rom_array[18902] = 32'hFFFFFFF0;
    // rom_array[18903] = 32'hFFFFFFF0;
    // rom_array[18904] = 32'hFFFFFFF0;
    // rom_array[18905] = 32'hFFFFFFF1;
    // rom_array[18906] = 32'hFFFFFFF1;
    // rom_array[18907] = 32'hFFFFFFF1;
    // rom_array[18908] = 32'hFFFFFFF1;
    // rom_array[18909] = 32'hFFFFFFF0;
    // rom_array[18910] = 32'hFFFFFFF0;
    // rom_array[18911] = 32'hFFFFFFF0;
    // rom_array[18912] = 32'hFFFFFFF0;
    // rom_array[18913] = 32'hFFFFFFF1;
    // rom_array[18914] = 32'hFFFFFFF1;
    // rom_array[18915] = 32'hFFFFFFF1;
    // rom_array[18916] = 32'hFFFFFFF1;
    // rom_array[18917] = 32'hFFFFFFF0;
    // rom_array[18918] = 32'hFFFFFFF0;
    // rom_array[18919] = 32'hFFFFFFF0;
    // rom_array[18920] = 32'hFFFFFFF0;
    // rom_array[18921] = 32'hFFFFFFF1;
    // rom_array[18922] = 32'hFFFFFFF1;
    // rom_array[18923] = 32'hFFFFFFF1;
    // rom_array[18924] = 32'hFFFFFFF1;
    // rom_array[18925] = 32'hFFFFFFF0;
    // rom_array[18926] = 32'hFFFFFFF0;
    // rom_array[18927] = 32'hFFFFFFF0;
    // rom_array[18928] = 32'hFFFFFFF0;
    // rom_array[18929] = 32'hFFFFFFF1;
    // rom_array[18930] = 32'hFFFFFFF1;
    // rom_array[18931] = 32'hFFFFFFF1;
    // rom_array[18932] = 32'hFFFFFFF1;
    // rom_array[18933] = 32'hFFFFFFF0;
    // rom_array[18934] = 32'hFFFFFFF0;
    // rom_array[18935] = 32'hFFFFFFF0;
    // rom_array[18936] = 32'hFFFFFFF0;
    // rom_array[18937] = 32'hFFFFFFF1;
    // rom_array[18938] = 32'hFFFFFFF1;
    // rom_array[18939] = 32'hFFFFFFF1;
    // rom_array[18940] = 32'hFFFFFFF1;
    // rom_array[18941] = 32'hFFFFFFF0;
    // rom_array[18942] = 32'hFFFFFFF0;
    // rom_array[18943] = 32'hFFFFFFF0;
    // rom_array[18944] = 32'hFFFFFFF0;
    // rom_array[18945] = 32'hFFFFFFF1;
    // rom_array[18946] = 32'hFFFFFFF1;
    // rom_array[18947] = 32'hFFFFFFF1;
    // rom_array[18948] = 32'hFFFFFFF1;
    // rom_array[18949] = 32'hFFFFFFF0;
    // rom_array[18950] = 32'hFFFFFFF0;
    // rom_array[18951] = 32'hFFFFFFF0;
    // rom_array[18952] = 32'hFFFFFFF0;
    // rom_array[18953] = 32'hFFFFFFF0;
    // rom_array[18954] = 32'hFFFFFFF0;
    // rom_array[18955] = 32'hFFFFFFF0;
    // rom_array[18956] = 32'hFFFFFFF0;
    // rom_array[18957] = 32'hFFFFFFF1;
    // rom_array[18958] = 32'hFFFFFFF1;
    // rom_array[18959] = 32'hFFFFFFF1;
    // rom_array[18960] = 32'hFFFFFFF1;
    // rom_array[18961] = 32'hFFFFFFF0;
    // rom_array[18962] = 32'hFFFFFFF0;
    // rom_array[18963] = 32'hFFFFFFF0;
    // rom_array[18964] = 32'hFFFFFFF0;
    // rom_array[18965] = 32'hFFFFFFF1;
    // rom_array[18966] = 32'hFFFFFFF1;
    // rom_array[18967] = 32'hFFFFFFF1;
    // rom_array[18968] = 32'hFFFFFFF1;
    // rom_array[18969] = 32'hFFFFFFF0;
    // rom_array[18970] = 32'hFFFFFFF0;
    // rom_array[18971] = 32'hFFFFFFF0;
    // rom_array[18972] = 32'hFFFFFFF0;
    // rom_array[18973] = 32'hFFFFFFF1;
    // rom_array[18974] = 32'hFFFFFFF1;
    // rom_array[18975] = 32'hFFFFFFF1;
    // rom_array[18976] = 32'hFFFFFFF1;
    // rom_array[18977] = 32'hFFFFFFF0;
    // rom_array[18978] = 32'hFFFFFFF0;
    // rom_array[18979] = 32'hFFFFFFF0;
    // rom_array[18980] = 32'hFFFFFFF0;
    // rom_array[18981] = 32'hFFFFFFF1;
    // rom_array[18982] = 32'hFFFFFFF1;
    // rom_array[18983] = 32'hFFFFFFF1;
    // rom_array[18984] = 32'hFFFFFFF1;
    // rom_array[18985] = 32'hFFFFFFF0;
    // rom_array[18986] = 32'hFFFFFFF0;
    // rom_array[18987] = 32'hFFFFFFF0;
    // rom_array[18988] = 32'hFFFFFFF0;
    // rom_array[18989] = 32'hFFFFFFF1;
    // rom_array[18990] = 32'hFFFFFFF1;
    // rom_array[18991] = 32'hFFFFFFF1;
    // rom_array[18992] = 32'hFFFFFFF1;
    // rom_array[18993] = 32'hFFFFFFF0;
    // rom_array[18994] = 32'hFFFFFFF0;
    // rom_array[18995] = 32'hFFFFFFF0;
    // rom_array[18996] = 32'hFFFFFFF0;
    // rom_array[18997] = 32'hFFFFFFF1;
    // rom_array[18998] = 32'hFFFFFFF1;
    // rom_array[18999] = 32'hFFFFFFF1;
    // rom_array[19000] = 32'hFFFFFFF1;
    // rom_array[19001] = 32'hFFFFFFF1;
    // rom_array[19002] = 32'hFFFFFFF1;
    // rom_array[19003] = 32'hFFFFFFF1;
    // rom_array[19004] = 32'hFFFFFFF1;
    // rom_array[19005] = 32'hFFFFFFF1;
    // rom_array[19006] = 32'hFFFFFFF1;
    // rom_array[19007] = 32'hFFFFFFF1;
    // rom_array[19008] = 32'hFFFFFFF1;
    // rom_array[19009] = 32'hFFFFFFF1;
    // rom_array[19010] = 32'hFFFFFFF1;
    // rom_array[19011] = 32'hFFFFFFF1;
    // rom_array[19012] = 32'hFFFFFFF1;
    // rom_array[19013] = 32'hFFFFFFF1;
    // rom_array[19014] = 32'hFFFFFFF1;
    // rom_array[19015] = 32'hFFFFFFF1;
    // rom_array[19016] = 32'hFFFFFFF1;
    // rom_array[19017] = 32'hFFFFFFF1;
    // rom_array[19018] = 32'hFFFFFFF1;
    // rom_array[19019] = 32'hFFFFFFF1;
    // rom_array[19020] = 32'hFFFFFFF1;
    // rom_array[19021] = 32'hFFFFFFF1;
    // rom_array[19022] = 32'hFFFFFFF1;
    // rom_array[19023] = 32'hFFFFFFF1;
    // rom_array[19024] = 32'hFFFFFFF1;
    // rom_array[19025] = 32'hFFFFFFF1;
    // rom_array[19026] = 32'hFFFFFFF1;
    // rom_array[19027] = 32'hFFFFFFF1;
    // rom_array[19028] = 32'hFFFFFFF1;
    // rom_array[19029] = 32'hFFFFFFF1;
    // rom_array[19030] = 32'hFFFFFFF1;
    // rom_array[19031] = 32'hFFFFFFF1;
    // rom_array[19032] = 32'hFFFFFFF1;
    // rom_array[19033] = 32'hFFFFFFF1;
    // rom_array[19034] = 32'hFFFFFFF1;
    // rom_array[19035] = 32'hFFFFFFF1;
    // rom_array[19036] = 32'hFFFFFFF1;
    // rom_array[19037] = 32'hFFFFFFF1;
    // rom_array[19038] = 32'hFFFFFFF1;
    // rom_array[19039] = 32'hFFFFFFF1;
    // rom_array[19040] = 32'hFFFFFFF1;
    // rom_array[19041] = 32'hFFFFFFF1;
    // rom_array[19042] = 32'hFFFFFFF1;
    // rom_array[19043] = 32'hFFFFFFF1;
    // rom_array[19044] = 32'hFFFFFFF1;
    // rom_array[19045] = 32'hFFFFFFF1;
    // rom_array[19046] = 32'hFFFFFFF1;
    // rom_array[19047] = 32'hFFFFFFF1;
    // rom_array[19048] = 32'hFFFFFFF1;
    // rom_array[19049] = 32'hFFFFFFF1;
    // rom_array[19050] = 32'hFFFFFFF1;
    // rom_array[19051] = 32'hFFFFFFF1;
    // rom_array[19052] = 32'hFFFFFFF1;
    // rom_array[19053] = 32'hFFFFFFF1;
    // rom_array[19054] = 32'hFFFFFFF1;
    // rom_array[19055] = 32'hFFFFFFF1;
    // rom_array[19056] = 32'hFFFFFFF1;
    // rom_array[19057] = 32'hFFFFFFF1;
    // rom_array[19058] = 32'hFFFFFFF1;
    // rom_array[19059] = 32'hFFFFFFF1;
    // rom_array[19060] = 32'hFFFFFFF1;
    // rom_array[19061] = 32'hFFFFFFF1;
    // rom_array[19062] = 32'hFFFFFFF1;
    // rom_array[19063] = 32'hFFFFFFF1;
    // rom_array[19064] = 32'hFFFFFFF1;
    // rom_array[19065] = 32'hFFFFFFF0;
    // rom_array[19066] = 32'hFFFFFFF0;
    // rom_array[19067] = 32'hFFFFFFF0;
    // rom_array[19068] = 32'hFFFFFFF0;
    // rom_array[19069] = 32'hFFFFFFF1;
    // rom_array[19070] = 32'hFFFFFFF1;
    // rom_array[19071] = 32'hFFFFFFF1;
    // rom_array[19072] = 32'hFFFFFFF1;
    // rom_array[19073] = 32'hFFFFFFF0;
    // rom_array[19074] = 32'hFFFFFFF0;
    // rom_array[19075] = 32'hFFFFFFF0;
    // rom_array[19076] = 32'hFFFFFFF0;
    // rom_array[19077] = 32'hFFFFFFF1;
    // rom_array[19078] = 32'hFFFFFFF1;
    // rom_array[19079] = 32'hFFFFFFF1;
    // rom_array[19080] = 32'hFFFFFFF1;
    // rom_array[19081] = 32'hFFFFFFF0;
    // rom_array[19082] = 32'hFFFFFFF0;
    // rom_array[19083] = 32'hFFFFFFF0;
    // rom_array[19084] = 32'hFFFFFFF0;
    // rom_array[19085] = 32'hFFFFFFF1;
    // rom_array[19086] = 32'hFFFFFFF1;
    // rom_array[19087] = 32'hFFFFFFF1;
    // rom_array[19088] = 32'hFFFFFFF1;
    // rom_array[19089] = 32'hFFFFFFF0;
    // rom_array[19090] = 32'hFFFFFFF0;
    // rom_array[19091] = 32'hFFFFFFF0;
    // rom_array[19092] = 32'hFFFFFFF0;
    // rom_array[19093] = 32'hFFFFFFF1;
    // rom_array[19094] = 32'hFFFFFFF1;
    // rom_array[19095] = 32'hFFFFFFF1;
    // rom_array[19096] = 32'hFFFFFFF1;
    // rom_array[19097] = 32'hFFFFFFF0;
    // rom_array[19098] = 32'hFFFFFFF0;
    // rom_array[19099] = 32'hFFFFFFF0;
    // rom_array[19100] = 32'hFFFFFFF0;
    // rom_array[19101] = 32'hFFFFFFF1;
    // rom_array[19102] = 32'hFFFFFFF1;
    // rom_array[19103] = 32'hFFFFFFF1;
    // rom_array[19104] = 32'hFFFFFFF1;
    // rom_array[19105] = 32'hFFFFFFF0;
    // rom_array[19106] = 32'hFFFFFFF0;
    // rom_array[19107] = 32'hFFFFFFF0;
    // rom_array[19108] = 32'hFFFFFFF0;
    // rom_array[19109] = 32'hFFFFFFF1;
    // rom_array[19110] = 32'hFFFFFFF1;
    // rom_array[19111] = 32'hFFFFFFF1;
    // rom_array[19112] = 32'hFFFFFFF1;
    // rom_array[19113] = 32'hFFFFFFF0;
    // rom_array[19114] = 32'hFFFFFFF0;
    // rom_array[19115] = 32'hFFFFFFF0;
    // rom_array[19116] = 32'hFFFFFFF0;
    // rom_array[19117] = 32'hFFFFFFF1;
    // rom_array[19118] = 32'hFFFFFFF1;
    // rom_array[19119] = 32'hFFFFFFF1;
    // rom_array[19120] = 32'hFFFFFFF1;
    // rom_array[19121] = 32'hFFFFFFF0;
    // rom_array[19122] = 32'hFFFFFFF0;
    // rom_array[19123] = 32'hFFFFFFF0;
    // rom_array[19124] = 32'hFFFFFFF0;
    // rom_array[19125] = 32'hFFFFFFF1;
    // rom_array[19126] = 32'hFFFFFFF1;
    // rom_array[19127] = 32'hFFFFFFF1;
    // rom_array[19128] = 32'hFFFFFFF1;
    // rom_array[19129] = 32'hFFFFFFF1;
    // rom_array[19130] = 32'hFFFFFFF1;
    // rom_array[19131] = 32'hFFFFFFF1;
    // rom_array[19132] = 32'hFFFFFFF1;
    // rom_array[19133] = 32'hFFFFFFF1;
    // rom_array[19134] = 32'hFFFFFFF1;
    // rom_array[19135] = 32'hFFFFFFF1;
    // rom_array[19136] = 32'hFFFFFFF1;
    // rom_array[19137] = 32'hFFFFFFF1;
    // rom_array[19138] = 32'hFFFFFFF1;
    // rom_array[19139] = 32'hFFFFFFF1;
    // rom_array[19140] = 32'hFFFFFFF1;
    // rom_array[19141] = 32'hFFFFFFF1;
    // rom_array[19142] = 32'hFFFFFFF1;
    // rom_array[19143] = 32'hFFFFFFF1;
    // rom_array[19144] = 32'hFFFFFFF1;
    // rom_array[19145] = 32'hFFFFFFF1;
    // rom_array[19146] = 32'hFFFFFFF1;
    // rom_array[19147] = 32'hFFFFFFF1;
    // rom_array[19148] = 32'hFFFFFFF1;
    // rom_array[19149] = 32'hFFFFFFF1;
    // rom_array[19150] = 32'hFFFFFFF1;
    // rom_array[19151] = 32'hFFFFFFF1;
    // rom_array[19152] = 32'hFFFFFFF1;
    // rom_array[19153] = 32'hFFFFFFF1;
    // rom_array[19154] = 32'hFFFFFFF1;
    // rom_array[19155] = 32'hFFFFFFF1;
    // rom_array[19156] = 32'hFFFFFFF1;
    // rom_array[19157] = 32'hFFFFFFF1;
    // rom_array[19158] = 32'hFFFFFFF1;
    // rom_array[19159] = 32'hFFFFFFF1;
    // rom_array[19160] = 32'hFFFFFFF1;
    // rom_array[19161] = 32'hFFFFFFF1;
    // rom_array[19162] = 32'hFFFFFFF1;
    // rom_array[19163] = 32'hFFFFFFF1;
    // rom_array[19164] = 32'hFFFFFFF1;
    // rom_array[19165] = 32'hFFFFFFF1;
    // rom_array[19166] = 32'hFFFFFFF1;
    // rom_array[19167] = 32'hFFFFFFF1;
    // rom_array[19168] = 32'hFFFFFFF1;
    // rom_array[19169] = 32'hFFFFFFF1;
    // rom_array[19170] = 32'hFFFFFFF1;
    // rom_array[19171] = 32'hFFFFFFF1;
    // rom_array[19172] = 32'hFFFFFFF1;
    // rom_array[19173] = 32'hFFFFFFF1;
    // rom_array[19174] = 32'hFFFFFFF1;
    // rom_array[19175] = 32'hFFFFFFF1;
    // rom_array[19176] = 32'hFFFFFFF1;
    // rom_array[19177] = 32'hFFFFFFF1;
    // rom_array[19178] = 32'hFFFFFFF1;
    // rom_array[19179] = 32'hFFFFFFF1;
    // rom_array[19180] = 32'hFFFFFFF1;
    // rom_array[19181] = 32'hFFFFFFF1;
    // rom_array[19182] = 32'hFFFFFFF1;
    // rom_array[19183] = 32'hFFFFFFF1;
    // rom_array[19184] = 32'hFFFFFFF1;
    // rom_array[19185] = 32'hFFFFFFF1;
    // rom_array[19186] = 32'hFFFFFFF1;
    // rom_array[19187] = 32'hFFFFFFF1;
    // rom_array[19188] = 32'hFFFFFFF1;
    // rom_array[19189] = 32'hFFFFFFF1;
    // rom_array[19190] = 32'hFFFFFFF1;
    // rom_array[19191] = 32'hFFFFFFF1;
    // rom_array[19192] = 32'hFFFFFFF1;
    // rom_array[19193] = 32'hFFFFFFF1;
    // rom_array[19194] = 32'hFFFFFFF1;
    // rom_array[19195] = 32'hFFFFFFF1;
    // rom_array[19196] = 32'hFFFFFFF1;
    // rom_array[19197] = 32'hFFFFFFF0;
    // rom_array[19198] = 32'hFFFFFFF0;
    // rom_array[19199] = 32'hFFFFFFF0;
    // rom_array[19200] = 32'hFFFFFFF0;
    // rom_array[19201] = 32'hFFFFFFF1;
    // rom_array[19202] = 32'hFFFFFFF1;
    // rom_array[19203] = 32'hFFFFFFF1;
    // rom_array[19204] = 32'hFFFFFFF1;
    // rom_array[19205] = 32'hFFFFFFF0;
    // rom_array[19206] = 32'hFFFFFFF0;
    // rom_array[19207] = 32'hFFFFFFF0;
    // rom_array[19208] = 32'hFFFFFFF0;
    // rom_array[19209] = 32'hFFFFFFF1;
    // rom_array[19210] = 32'hFFFFFFF1;
    // rom_array[19211] = 32'hFFFFFFF1;
    // rom_array[19212] = 32'hFFFFFFF1;
    // rom_array[19213] = 32'hFFFFFFF0;
    // rom_array[19214] = 32'hFFFFFFF0;
    // rom_array[19215] = 32'hFFFFFFF0;
    // rom_array[19216] = 32'hFFFFFFF0;
    // rom_array[19217] = 32'hFFFFFFF1;
    // rom_array[19218] = 32'hFFFFFFF1;
    // rom_array[19219] = 32'hFFFFFFF1;
    // rom_array[19220] = 32'hFFFFFFF1;
    // rom_array[19221] = 32'hFFFFFFF0;
    // rom_array[19222] = 32'hFFFFFFF0;
    // rom_array[19223] = 32'hFFFFFFF0;
    // rom_array[19224] = 32'hFFFFFFF0;
    // rom_array[19225] = 32'hFFFFFFF1;
    // rom_array[19226] = 32'hFFFFFFF1;
    // rom_array[19227] = 32'hFFFFFFF1;
    // rom_array[19228] = 32'hFFFFFFF1;
    // rom_array[19229] = 32'hFFFFFFF0;
    // rom_array[19230] = 32'hFFFFFFF0;
    // rom_array[19231] = 32'hFFFFFFF0;
    // rom_array[19232] = 32'hFFFFFFF0;
    // rom_array[19233] = 32'hFFFFFFF1;
    // rom_array[19234] = 32'hFFFFFFF1;
    // rom_array[19235] = 32'hFFFFFFF1;
    // rom_array[19236] = 32'hFFFFFFF1;
    // rom_array[19237] = 32'hFFFFFFF0;
    // rom_array[19238] = 32'hFFFFFFF0;
    // rom_array[19239] = 32'hFFFFFFF0;
    // rom_array[19240] = 32'hFFFFFFF0;
    // rom_array[19241] = 32'hFFFFFFF1;
    // rom_array[19242] = 32'hFFFFFFF1;
    // rom_array[19243] = 32'hFFFFFFF1;
    // rom_array[19244] = 32'hFFFFFFF1;
    // rom_array[19245] = 32'hFFFFFFF0;
    // rom_array[19246] = 32'hFFFFFFF0;
    // rom_array[19247] = 32'hFFFFFFF0;
    // rom_array[19248] = 32'hFFFFFFF0;
    // rom_array[19249] = 32'hFFFFFFF1;
    // rom_array[19250] = 32'hFFFFFFF1;
    // rom_array[19251] = 32'hFFFFFFF1;
    // rom_array[19252] = 32'hFFFFFFF1;
    // rom_array[19253] = 32'hFFFFFFF0;
    // rom_array[19254] = 32'hFFFFFFF0;
    // rom_array[19255] = 32'hFFFFFFF0;
    // rom_array[19256] = 32'hFFFFFFF0;
    // rom_array[19257] = 32'hFFFFFFF1;
    // rom_array[19258] = 32'hFFFFFFF1;
    // rom_array[19259] = 32'hFFFFFFF1;
    // rom_array[19260] = 32'hFFFFFFF1;
    // rom_array[19261] = 32'hFFFFFFF0;
    // rom_array[19262] = 32'hFFFFFFF0;
    // rom_array[19263] = 32'hFFFFFFF0;
    // rom_array[19264] = 32'hFFFFFFF0;
    // rom_array[19265] = 32'hFFFFFFF1;
    // rom_array[19266] = 32'hFFFFFFF1;
    // rom_array[19267] = 32'hFFFFFFF1;
    // rom_array[19268] = 32'hFFFFFFF1;
    // rom_array[19269] = 32'hFFFFFFF0;
    // rom_array[19270] = 32'hFFFFFFF0;
    // rom_array[19271] = 32'hFFFFFFF0;
    // rom_array[19272] = 32'hFFFFFFF0;
    // rom_array[19273] = 32'hFFFFFFF1;
    // rom_array[19274] = 32'hFFFFFFF1;
    // rom_array[19275] = 32'hFFFFFFF1;
    // rom_array[19276] = 32'hFFFFFFF1;
    // rom_array[19277] = 32'hFFFFFFF0;
    // rom_array[19278] = 32'hFFFFFFF0;
    // rom_array[19279] = 32'hFFFFFFF0;
    // rom_array[19280] = 32'hFFFFFFF0;
    // rom_array[19281] = 32'hFFFFFFF1;
    // rom_array[19282] = 32'hFFFFFFF1;
    // rom_array[19283] = 32'hFFFFFFF1;
    // rom_array[19284] = 32'hFFFFFFF1;
    // rom_array[19285] = 32'hFFFFFFF0;
    // rom_array[19286] = 32'hFFFFFFF0;
    // rom_array[19287] = 32'hFFFFFFF0;
    // rom_array[19288] = 32'hFFFFFFF0;
    // rom_array[19289] = 32'hFFFFFFF1;
    // rom_array[19290] = 32'hFFFFFFF1;
    // rom_array[19291] = 32'hFFFFFFF1;
    // rom_array[19292] = 32'hFFFFFFF1;
    // rom_array[19293] = 32'hFFFFFFF0;
    // rom_array[19294] = 32'hFFFFFFF0;
    // rom_array[19295] = 32'hFFFFFFF0;
    // rom_array[19296] = 32'hFFFFFFF0;
    // rom_array[19297] = 32'hFFFFFFF1;
    // rom_array[19298] = 32'hFFFFFFF1;
    // rom_array[19299] = 32'hFFFFFFF1;
    // rom_array[19300] = 32'hFFFFFFF1;
    // rom_array[19301] = 32'hFFFFFFF0;
    // rom_array[19302] = 32'hFFFFFFF0;
    // rom_array[19303] = 32'hFFFFFFF0;
    // rom_array[19304] = 32'hFFFFFFF0;
    // rom_array[19305] = 32'hFFFFFFF1;
    // rom_array[19306] = 32'hFFFFFFF1;
    // rom_array[19307] = 32'hFFFFFFF1;
    // rom_array[19308] = 32'hFFFFFFF1;
    // rom_array[19309] = 32'hFFFFFFF0;
    // rom_array[19310] = 32'hFFFFFFF0;
    // rom_array[19311] = 32'hFFFFFFF0;
    // rom_array[19312] = 32'hFFFFFFF0;
    // rom_array[19313] = 32'hFFFFFFF1;
    // rom_array[19314] = 32'hFFFFFFF1;
    // rom_array[19315] = 32'hFFFFFFF1;
    // rom_array[19316] = 32'hFFFFFFF1;
    // rom_array[19317] = 32'hFFFFFFF0;
    // rom_array[19318] = 32'hFFFFFFF0;
    // rom_array[19319] = 32'hFFFFFFF0;
    // rom_array[19320] = 32'hFFFFFFF0;
    // rom_array[19321] = 32'hFFFFFFF0;
    // rom_array[19322] = 32'hFFFFFFF0;
    // rom_array[19323] = 32'hFFFFFFF0;
    // rom_array[19324] = 32'hFFFFFFF0;
    // rom_array[19325] = 32'hFFFFFFF0;
    // rom_array[19326] = 32'hFFFFFFF0;
    // rom_array[19327] = 32'hFFFFFFF1;
    // rom_array[19328] = 32'hFFFFFFF1;
    // rom_array[19329] = 32'hFFFFFFF0;
    // rom_array[19330] = 32'hFFFFFFF0;
    // rom_array[19331] = 32'hFFFFFFF0;
    // rom_array[19332] = 32'hFFFFFFF0;
    // rom_array[19333] = 32'hFFFFFFF0;
    // rom_array[19334] = 32'hFFFFFFF0;
    // rom_array[19335] = 32'hFFFFFFF1;
    // rom_array[19336] = 32'hFFFFFFF1;
    // rom_array[19337] = 32'hFFFFFFF0;
    // rom_array[19338] = 32'hFFFFFFF0;
    // rom_array[19339] = 32'hFFFFFFF0;
    // rom_array[19340] = 32'hFFFFFFF0;
    // rom_array[19341] = 32'hFFFFFFF1;
    // rom_array[19342] = 32'hFFFFFFF1;
    // rom_array[19343] = 32'hFFFFFFF1;
    // rom_array[19344] = 32'hFFFFFFF1;
    // rom_array[19345] = 32'hFFFFFFF0;
    // rom_array[19346] = 32'hFFFFFFF0;
    // rom_array[19347] = 32'hFFFFFFF0;
    // rom_array[19348] = 32'hFFFFFFF0;
    // rom_array[19349] = 32'hFFFFFFF1;
    // rom_array[19350] = 32'hFFFFFFF1;
    // rom_array[19351] = 32'hFFFFFFF1;
    // rom_array[19352] = 32'hFFFFFFF1;
    // rom_array[19353] = 32'hFFFFFFF0;
    // rom_array[19354] = 32'hFFFFFFF0;
    // rom_array[19355] = 32'hFFFFFFF1;
    // rom_array[19356] = 32'hFFFFFFF1;
    // rom_array[19357] = 32'hFFFFFFF0;
    // rom_array[19358] = 32'hFFFFFFF0;
    // rom_array[19359] = 32'hFFFFFFF1;
    // rom_array[19360] = 32'hFFFFFFF1;
    // rom_array[19361] = 32'hFFFFFFF0;
    // rom_array[19362] = 32'hFFFFFFF0;
    // rom_array[19363] = 32'hFFFFFFF1;
    // rom_array[19364] = 32'hFFFFFFF1;
    // rom_array[19365] = 32'hFFFFFFF0;
    // rom_array[19366] = 32'hFFFFFFF0;
    // rom_array[19367] = 32'hFFFFFFF1;
    // rom_array[19368] = 32'hFFFFFFF1;
    // rom_array[19369] = 32'hFFFFFFF0;
    // rom_array[19370] = 32'hFFFFFFF0;
    // rom_array[19371] = 32'hFFFFFFF0;
    // rom_array[19372] = 32'hFFFFFFF0;
    // rom_array[19373] = 32'hFFFFFFF1;
    // rom_array[19374] = 32'hFFFFFFF1;
    // rom_array[19375] = 32'hFFFFFFF1;
    // rom_array[19376] = 32'hFFFFFFF1;
    // rom_array[19377] = 32'hFFFFFFF0;
    // rom_array[19378] = 32'hFFFFFFF0;
    // rom_array[19379] = 32'hFFFFFFF0;
    // rom_array[19380] = 32'hFFFFFFF0;
    // rom_array[19381] = 32'hFFFFFFF1;
    // rom_array[19382] = 32'hFFFFFFF1;
    // rom_array[19383] = 32'hFFFFFFF1;
    // rom_array[19384] = 32'hFFFFFFF1;
    // rom_array[19385] = 32'hFFFFFFF0;
    // rom_array[19386] = 32'hFFFFFFF0;
    // rom_array[19387] = 32'hFFFFFFF0;
    // rom_array[19388] = 32'hFFFFFFF0;
    // rom_array[19389] = 32'hFFFFFFF1;
    // rom_array[19390] = 32'hFFFFFFF1;
    // rom_array[19391] = 32'hFFFFFFF1;
    // rom_array[19392] = 32'hFFFFFFF1;
    // rom_array[19393] = 32'hFFFFFFF0;
    // rom_array[19394] = 32'hFFFFFFF0;
    // rom_array[19395] = 32'hFFFFFFF0;
    // rom_array[19396] = 32'hFFFFFFF0;
    // rom_array[19397] = 32'hFFFFFFF1;
    // rom_array[19398] = 32'hFFFFFFF1;
    // rom_array[19399] = 32'hFFFFFFF1;
    // rom_array[19400] = 32'hFFFFFFF1;
    // rom_array[19401] = 32'hFFFFFFF0;
    // rom_array[19402] = 32'hFFFFFFF0;
    // rom_array[19403] = 32'hFFFFFFF1;
    // rom_array[19404] = 32'hFFFFFFF1;
    // rom_array[19405] = 32'hFFFFFFF0;
    // rom_array[19406] = 32'hFFFFFFF0;
    // rom_array[19407] = 32'hFFFFFFF1;
    // rom_array[19408] = 32'hFFFFFFF1;
    // rom_array[19409] = 32'hFFFFFFF0;
    // rom_array[19410] = 32'hFFFFFFF0;
    // rom_array[19411] = 32'hFFFFFFF1;
    // rom_array[19412] = 32'hFFFFFFF1;
    // rom_array[19413] = 32'hFFFFFFF0;
    // rom_array[19414] = 32'hFFFFFFF0;
    // rom_array[19415] = 32'hFFFFFFF1;
    // rom_array[19416] = 32'hFFFFFFF1;
    // rom_array[19417] = 32'hFFFFFFF0;
    // rom_array[19418] = 32'hFFFFFFF0;
    // rom_array[19419] = 32'hFFFFFFF1;
    // rom_array[19420] = 32'hFFFFFFF1;
    // rom_array[19421] = 32'hFFFFFFF0;
    // rom_array[19422] = 32'hFFFFFFF0;
    // rom_array[19423] = 32'hFFFFFFF1;
    // rom_array[19424] = 32'hFFFFFFF1;
    // rom_array[19425] = 32'hFFFFFFF0;
    // rom_array[19426] = 32'hFFFFFFF0;
    // rom_array[19427] = 32'hFFFFFFF1;
    // rom_array[19428] = 32'hFFFFFFF1;
    // rom_array[19429] = 32'hFFFFFFF0;
    // rom_array[19430] = 32'hFFFFFFF0;
    // rom_array[19431] = 32'hFFFFFFF1;
    // rom_array[19432] = 32'hFFFFFFF1;
    // rom_array[19433] = 32'hFFFFFFF0;
    // rom_array[19434] = 32'hFFFFFFF0;
    // rom_array[19435] = 32'hFFFFFFF1;
    // rom_array[19436] = 32'hFFFFFFF1;
    // rom_array[19437] = 32'hFFFFFFF0;
    // rom_array[19438] = 32'hFFFFFFF0;
    // rom_array[19439] = 32'hFFFFFFF0;
    // rom_array[19440] = 32'hFFFFFFF0;
    // rom_array[19441] = 32'hFFFFFFF0;
    // rom_array[19442] = 32'hFFFFFFF0;
    // rom_array[19443] = 32'hFFFFFFF1;
    // rom_array[19444] = 32'hFFFFFFF1;
    // rom_array[19445] = 32'hFFFFFFF0;
    // rom_array[19446] = 32'hFFFFFFF0;
    // rom_array[19447] = 32'hFFFFFFF0;
    // rom_array[19448] = 32'hFFFFFFF0;
    // rom_array[19449] = 32'hFFFFFFF1;
    // rom_array[19450] = 32'hFFFFFFF1;
    // rom_array[19451] = 32'hFFFFFFF1;
    // rom_array[19452] = 32'hFFFFFFF1;
    // rom_array[19453] = 32'hFFFFFFF0;
    // rom_array[19454] = 32'hFFFFFFF0;
    // rom_array[19455] = 32'hFFFFFFF0;
    // rom_array[19456] = 32'hFFFFFFF0;
    // rom_array[19457] = 32'hFFFFFFF1;
    // rom_array[19458] = 32'hFFFFFFF1;
    // rom_array[19459] = 32'hFFFFFFF1;
    // rom_array[19460] = 32'hFFFFFFF1;
    // rom_array[19461] = 32'hFFFFFFF0;
    // rom_array[19462] = 32'hFFFFFFF0;
    // rom_array[19463] = 32'hFFFFFFF0;
    // rom_array[19464] = 32'hFFFFFFF0;
    // rom_array[19465] = 32'hFFFFFFF1;
    // rom_array[19466] = 32'hFFFFFFF1;
    // rom_array[19467] = 32'hFFFFFFF1;
    // rom_array[19468] = 32'hFFFFFFF1;
    // rom_array[19469] = 32'hFFFFFFF0;
    // rom_array[19470] = 32'hFFFFFFF0;
    // rom_array[19471] = 32'hFFFFFFF0;
    // rom_array[19472] = 32'hFFFFFFF0;
    // rom_array[19473] = 32'hFFFFFFF1;
    // rom_array[19474] = 32'hFFFFFFF1;
    // rom_array[19475] = 32'hFFFFFFF1;
    // rom_array[19476] = 32'hFFFFFFF1;
    // rom_array[19477] = 32'hFFFFFFF0;
    // rom_array[19478] = 32'hFFFFFFF0;
    // rom_array[19479] = 32'hFFFFFFF0;
    // rom_array[19480] = 32'hFFFFFFF0;
    // rom_array[19481] = 32'hFFFFFFF1;
    // rom_array[19482] = 32'hFFFFFFF1;
    // rom_array[19483] = 32'hFFFFFFF1;
    // rom_array[19484] = 32'hFFFFFFF1;
    // rom_array[19485] = 32'hFFFFFFF0;
    // rom_array[19486] = 32'hFFFFFFF0;
    // rom_array[19487] = 32'hFFFFFFF0;
    // rom_array[19488] = 32'hFFFFFFF0;
    // rom_array[19489] = 32'hFFFFFFF1;
    // rom_array[19490] = 32'hFFFFFFF1;
    // rom_array[19491] = 32'hFFFFFFF1;
    // rom_array[19492] = 32'hFFFFFFF1;
    // rom_array[19493] = 32'hFFFFFFF0;
    // rom_array[19494] = 32'hFFFFFFF0;
    // rom_array[19495] = 32'hFFFFFFF0;
    // rom_array[19496] = 32'hFFFFFFF0;
    // rom_array[19497] = 32'hFFFFFFF0;
    // rom_array[19498] = 32'hFFFFFFF0;
    // rom_array[19499] = 32'hFFFFFFF0;
    // rom_array[19500] = 32'hFFFFFFF0;
    // rom_array[19501] = 32'hFFFFFFF1;
    // rom_array[19502] = 32'hFFFFFFF1;
    // rom_array[19503] = 32'hFFFFFFF1;
    // rom_array[19504] = 32'hFFFFFFF1;
    // rom_array[19505] = 32'hFFFFFFF0;
    // rom_array[19506] = 32'hFFFFFFF0;
    // rom_array[19507] = 32'hFFFFFFF0;
    // rom_array[19508] = 32'hFFFFFFF0;
    // rom_array[19509] = 32'hFFFFFFF1;
    // rom_array[19510] = 32'hFFFFFFF1;
    // rom_array[19511] = 32'hFFFFFFF1;
    // rom_array[19512] = 32'hFFFFFFF1;
    // rom_array[19513] = 32'hFFFFFFF0;
    // rom_array[19514] = 32'hFFFFFFF0;
    // rom_array[19515] = 32'hFFFFFFF0;
    // rom_array[19516] = 32'hFFFFFFF0;
    // rom_array[19517] = 32'hFFFFFFF1;
    // rom_array[19518] = 32'hFFFFFFF1;
    // rom_array[19519] = 32'hFFFFFFF1;
    // rom_array[19520] = 32'hFFFFFFF1;
    // rom_array[19521] = 32'hFFFFFFF0;
    // rom_array[19522] = 32'hFFFFFFF0;
    // rom_array[19523] = 32'hFFFFFFF0;
    // rom_array[19524] = 32'hFFFFFFF0;
    // rom_array[19525] = 32'hFFFFFFF1;
    // rom_array[19526] = 32'hFFFFFFF1;
    // rom_array[19527] = 32'hFFFFFFF1;
    // rom_array[19528] = 32'hFFFFFFF1;
    // rom_array[19529] = 32'hFFFFFFF0;
    // rom_array[19530] = 32'hFFFFFFF0;
    // rom_array[19531] = 32'hFFFFFFF0;
    // rom_array[19532] = 32'hFFFFFFF0;
    // rom_array[19533] = 32'hFFFFFFF1;
    // rom_array[19534] = 32'hFFFFFFF1;
    // rom_array[19535] = 32'hFFFFFFF1;
    // rom_array[19536] = 32'hFFFFFFF1;
    // rom_array[19537] = 32'hFFFFFFF0;
    // rom_array[19538] = 32'hFFFFFFF0;
    // rom_array[19539] = 32'hFFFFFFF0;
    // rom_array[19540] = 32'hFFFFFFF0;
    // rom_array[19541] = 32'hFFFFFFF1;
    // rom_array[19542] = 32'hFFFFFFF1;
    // rom_array[19543] = 32'hFFFFFFF1;
    // rom_array[19544] = 32'hFFFFFFF1;
    // rom_array[19545] = 32'hFFFFFFF0;
    // rom_array[19546] = 32'hFFFFFFF0;
    // rom_array[19547] = 32'hFFFFFFF0;
    // rom_array[19548] = 32'hFFFFFFF0;
    // rom_array[19549] = 32'hFFFFFFF1;
    // rom_array[19550] = 32'hFFFFFFF1;
    // rom_array[19551] = 32'hFFFFFFF1;
    // rom_array[19552] = 32'hFFFFFFF1;
    // rom_array[19553] = 32'hFFFFFFF0;
    // rom_array[19554] = 32'hFFFFFFF0;
    // rom_array[19555] = 32'hFFFFFFF0;
    // rom_array[19556] = 32'hFFFFFFF0;
    // rom_array[19557] = 32'hFFFFFFF1;
    // rom_array[19558] = 32'hFFFFFFF1;
    // rom_array[19559] = 32'hFFFFFFF1;
    // rom_array[19560] = 32'hFFFFFFF1;
    // rom_array[19561] = 32'hFFFFFFF0;
    // rom_array[19562] = 32'hFFFFFFF0;
    // rom_array[19563] = 32'hFFFFFFF0;
    // rom_array[19564] = 32'hFFFFFFF0;
    // rom_array[19565] = 32'hFFFFFFF1;
    // rom_array[19566] = 32'hFFFFFFF1;
    // rom_array[19567] = 32'hFFFFFFF1;
    // rom_array[19568] = 32'hFFFFFFF1;
    // rom_array[19569] = 32'hFFFFFFF0;
    // rom_array[19570] = 32'hFFFFFFF0;
    // rom_array[19571] = 32'hFFFFFFF0;
    // rom_array[19572] = 32'hFFFFFFF0;
    // rom_array[19573] = 32'hFFFFFFF1;
    // rom_array[19574] = 32'hFFFFFFF1;
    // rom_array[19575] = 32'hFFFFFFF1;
    // rom_array[19576] = 32'hFFFFFFF1;
    // rom_array[19577] = 32'hFFFFFFF0;
    // rom_array[19578] = 32'hFFFFFFF0;
    // rom_array[19579] = 32'hFFFFFFF0;
    // rom_array[19580] = 32'hFFFFFFF0;
    // rom_array[19581] = 32'hFFFFFFF1;
    // rom_array[19582] = 32'hFFFFFFF1;
    // rom_array[19583] = 32'hFFFFFFF1;
    // rom_array[19584] = 32'hFFFFFFF1;
    // rom_array[19585] = 32'hFFFFFFF0;
    // rom_array[19586] = 32'hFFFFFFF0;
    // rom_array[19587] = 32'hFFFFFFF0;
    // rom_array[19588] = 32'hFFFFFFF0;
    // rom_array[19589] = 32'hFFFFFFF1;
    // rom_array[19590] = 32'hFFFFFFF1;
    // rom_array[19591] = 32'hFFFFFFF1;
    // rom_array[19592] = 32'hFFFFFFF1;
    // rom_array[19593] = 32'hFFFFFFF0;
    // rom_array[19594] = 32'hFFFFFFF0;
    // rom_array[19595] = 32'hFFFFFFF0;
    // rom_array[19596] = 32'hFFFFFFF0;
    // rom_array[19597] = 32'hFFFFFFF1;
    // rom_array[19598] = 32'hFFFFFFF1;
    // rom_array[19599] = 32'hFFFFFFF1;
    // rom_array[19600] = 32'hFFFFFFF1;
    // rom_array[19601] = 32'hFFFFFFF0;
    // rom_array[19602] = 32'hFFFFFFF0;
    // rom_array[19603] = 32'hFFFFFFF0;
    // rom_array[19604] = 32'hFFFFFFF0;
    // rom_array[19605] = 32'hFFFFFFF1;
    // rom_array[19606] = 32'hFFFFFFF1;
    // rom_array[19607] = 32'hFFFFFFF1;
    // rom_array[19608] = 32'hFFFFFFF1;
    // rom_array[19609] = 32'hFFFFFFF0;
    // rom_array[19610] = 32'hFFFFFFF0;
    // rom_array[19611] = 32'hFFFFFFF0;
    // rom_array[19612] = 32'hFFFFFFF0;
    // rom_array[19613] = 32'hFFFFFFF1;
    // rom_array[19614] = 32'hFFFFFFF1;
    // rom_array[19615] = 32'hFFFFFFF1;
    // rom_array[19616] = 32'hFFFFFFF1;
    // rom_array[19617] = 32'hFFFFFFF0;
    // rom_array[19618] = 32'hFFFFFFF0;
    // rom_array[19619] = 32'hFFFFFFF0;
    // rom_array[19620] = 32'hFFFFFFF0;
    // rom_array[19621] = 32'hFFFFFFF1;
    // rom_array[19622] = 32'hFFFFFFF1;
    // rom_array[19623] = 32'hFFFFFFF1;
    // rom_array[19624] = 32'hFFFFFFF1;
    // rom_array[19625] = 32'hFFFFFFF1;
    // rom_array[19626] = 32'hFFFFFFF1;
    // rom_array[19627] = 32'hFFFFFFF1;
    // rom_array[19628] = 32'hFFFFFFF1;
    // rom_array[19629] = 32'hFFFFFFF0;
    // rom_array[19630] = 32'hFFFFFFF0;
    // rom_array[19631] = 32'hFFFFFFF0;
    // rom_array[19632] = 32'hFFFFFFF0;
    // rom_array[19633] = 32'hFFFFFFF1;
    // rom_array[19634] = 32'hFFFFFFF1;
    // rom_array[19635] = 32'hFFFFFFF1;
    // rom_array[19636] = 32'hFFFFFFF1;
    // rom_array[19637] = 32'hFFFFFFF0;
    // rom_array[19638] = 32'hFFFFFFF0;
    // rom_array[19639] = 32'hFFFFFFF0;
    // rom_array[19640] = 32'hFFFFFFF0;
    // rom_array[19641] = 32'hFFFFFFF1;
    // rom_array[19642] = 32'hFFFFFFF1;
    // rom_array[19643] = 32'hFFFFFFF1;
    // rom_array[19644] = 32'hFFFFFFF1;
    // rom_array[19645] = 32'hFFFFFFF0;
    // rom_array[19646] = 32'hFFFFFFF0;
    // rom_array[19647] = 32'hFFFFFFF0;
    // rom_array[19648] = 32'hFFFFFFF0;
    // rom_array[19649] = 32'hFFFFFFF1;
    // rom_array[19650] = 32'hFFFFFFF1;
    // rom_array[19651] = 32'hFFFFFFF1;
    // rom_array[19652] = 32'hFFFFFFF1;
    // rom_array[19653] = 32'hFFFFFFF0;
    // rom_array[19654] = 32'hFFFFFFF0;
    // rom_array[19655] = 32'hFFFFFFF0;
    // rom_array[19656] = 32'hFFFFFFF0;
    // rom_array[19657] = 32'hFFFFFFF1;
    // rom_array[19658] = 32'hFFFFFFF1;
    // rom_array[19659] = 32'hFFFFFFF1;
    // rom_array[19660] = 32'hFFFFFFF1;
    // rom_array[19661] = 32'hFFFFFFF0;
    // rom_array[19662] = 32'hFFFFFFF0;
    // rom_array[19663] = 32'hFFFFFFF0;
    // rom_array[19664] = 32'hFFFFFFF0;
    // rom_array[19665] = 32'hFFFFFFF1;
    // rom_array[19666] = 32'hFFFFFFF1;
    // rom_array[19667] = 32'hFFFFFFF1;
    // rom_array[19668] = 32'hFFFFFFF1;
    // rom_array[19669] = 32'hFFFFFFF0;
    // rom_array[19670] = 32'hFFFFFFF0;
    // rom_array[19671] = 32'hFFFFFFF0;
    // rom_array[19672] = 32'hFFFFFFF0;
    // rom_array[19673] = 32'hFFFFFFF1;
    // rom_array[19674] = 32'hFFFFFFF1;
    // rom_array[19675] = 32'hFFFFFFF1;
    // rom_array[19676] = 32'hFFFFFFF1;
    // rom_array[19677] = 32'hFFFFFFF0;
    // rom_array[19678] = 32'hFFFFFFF0;
    // rom_array[19679] = 32'hFFFFFFF0;
    // rom_array[19680] = 32'hFFFFFFF0;
    // rom_array[19681] = 32'hFFFFFFF1;
    // rom_array[19682] = 32'hFFFFFFF1;
    // rom_array[19683] = 32'hFFFFFFF1;
    // rom_array[19684] = 32'hFFFFFFF1;
    // rom_array[19685] = 32'hFFFFFFF0;
    // rom_array[19686] = 32'hFFFFFFF0;
    // rom_array[19687] = 32'hFFFFFFF0;
    // rom_array[19688] = 32'hFFFFFFF0;
    // rom_array[19689] = 32'hFFFFFFF1;
    // rom_array[19690] = 32'hFFFFFFF1;
    // rom_array[19691] = 32'hFFFFFFF1;
    // rom_array[19692] = 32'hFFFFFFF1;
    // rom_array[19693] = 32'hFFFFFFF0;
    // rom_array[19694] = 32'hFFFFFFF0;
    // rom_array[19695] = 32'hFFFFFFF1;
    // rom_array[19696] = 32'hFFFFFFF1;
    // rom_array[19697] = 32'hFFFFFFF1;
    // rom_array[19698] = 32'hFFFFFFF1;
    // rom_array[19699] = 32'hFFFFFFF1;
    // rom_array[19700] = 32'hFFFFFFF1;
    // rom_array[19701] = 32'hFFFFFFF0;
    // rom_array[19702] = 32'hFFFFFFF0;
    // rom_array[19703] = 32'hFFFFFFF1;
    // rom_array[19704] = 32'hFFFFFFF1;
    // rom_array[19705] = 32'hFFFFFFF1;
    // rom_array[19706] = 32'hFFFFFFF1;
    // rom_array[19707] = 32'hFFFFFFF1;
    // rom_array[19708] = 32'hFFFFFFF1;
    // rom_array[19709] = 32'hFFFFFFF1;
    // rom_array[19710] = 32'hFFFFFFF1;
    // rom_array[19711] = 32'hFFFFFFF1;
    // rom_array[19712] = 32'hFFFFFFF1;
    // rom_array[19713] = 32'hFFFFFFF1;
    // rom_array[19714] = 32'hFFFFFFF1;
    // rom_array[19715] = 32'hFFFFFFF1;
    // rom_array[19716] = 32'hFFFFFFF1;
    // rom_array[19717] = 32'hFFFFFFF1;
    // rom_array[19718] = 32'hFFFFFFF1;
    // rom_array[19719] = 32'hFFFFFFF1;
    // rom_array[19720] = 32'hFFFFFFF1;
    // rom_array[19721] = 32'hFFFFFFF0;
    // rom_array[19722] = 32'hFFFFFFF0;
    // rom_array[19723] = 32'hFFFFFFF1;
    // rom_array[19724] = 32'hFFFFFFF1;
    // rom_array[19725] = 32'hFFFFFFF0;
    // rom_array[19726] = 32'hFFFFFFF0;
    // rom_array[19727] = 32'hFFFFFFF1;
    // rom_array[19728] = 32'hFFFFFFF1;
    // rom_array[19729] = 32'hFFFFFFF0;
    // rom_array[19730] = 32'hFFFFFFF0;
    // rom_array[19731] = 32'hFFFFFFF1;
    // rom_array[19732] = 32'hFFFFFFF1;
    // rom_array[19733] = 32'hFFFFFFF0;
    // rom_array[19734] = 32'hFFFFFFF0;
    // rom_array[19735] = 32'hFFFFFFF1;
    // rom_array[19736] = 32'hFFFFFFF1;
    // rom_array[19737] = 32'hFFFFFFF1;
    // rom_array[19738] = 32'hFFFFFFF1;
    // rom_array[19739] = 32'hFFFFFFF1;
    // rom_array[19740] = 32'hFFFFFFF1;
    // rom_array[19741] = 32'hFFFFFFF1;
    // rom_array[19742] = 32'hFFFFFFF1;
    // rom_array[19743] = 32'hFFFFFFF1;
    // rom_array[19744] = 32'hFFFFFFF1;
    // rom_array[19745] = 32'hFFFFFFF1;
    // rom_array[19746] = 32'hFFFFFFF1;
    // rom_array[19747] = 32'hFFFFFFF1;
    // rom_array[19748] = 32'hFFFFFFF1;
    // rom_array[19749] = 32'hFFFFFFF1;
    // rom_array[19750] = 32'hFFFFFFF1;
    // rom_array[19751] = 32'hFFFFFFF1;
    // rom_array[19752] = 32'hFFFFFFF1;
    // rom_array[19753] = 32'hFFFFFFF1;
    // rom_array[19754] = 32'hFFFFFFF1;
    // rom_array[19755] = 32'hFFFFFFF1;
    // rom_array[19756] = 32'hFFFFFFF1;
    // rom_array[19757] = 32'hFFFFFFF1;
    // rom_array[19758] = 32'hFFFFFFF1;
    // rom_array[19759] = 32'hFFFFFFF1;
    // rom_array[19760] = 32'hFFFFFFF1;
    // rom_array[19761] = 32'hFFFFFFF1;
    // rom_array[19762] = 32'hFFFFFFF1;
    // rom_array[19763] = 32'hFFFFFFF1;
    // rom_array[19764] = 32'hFFFFFFF1;
    // rom_array[19765] = 32'hFFFFFFF1;
    // rom_array[19766] = 32'hFFFFFFF1;
    // rom_array[19767] = 32'hFFFFFFF1;
    // rom_array[19768] = 32'hFFFFFFF1;
    // rom_array[19769] = 32'hFFFFFFF0;
    // rom_array[19770] = 32'hFFFFFFF0;
    // rom_array[19771] = 32'hFFFFFFF1;
    // rom_array[19772] = 32'hFFFFFFF1;
    // rom_array[19773] = 32'hFFFFFFF0;
    // rom_array[19774] = 32'hFFFFFFF0;
    // rom_array[19775] = 32'hFFFFFFF1;
    // rom_array[19776] = 32'hFFFFFFF1;
    // rom_array[19777] = 32'hFFFFFFF0;
    // rom_array[19778] = 32'hFFFFFFF0;
    // rom_array[19779] = 32'hFFFFFFF1;
    // rom_array[19780] = 32'hFFFFFFF1;
    // rom_array[19781] = 32'hFFFFFFF0;
    // rom_array[19782] = 32'hFFFFFFF0;
    // rom_array[19783] = 32'hFFFFFFF1;
    // rom_array[19784] = 32'hFFFFFFF1;
    // rom_array[19785] = 32'hFFFFFFF0;
    // rom_array[19786] = 32'hFFFFFFF0;
    // rom_array[19787] = 32'hFFFFFFF1;
    // rom_array[19788] = 32'hFFFFFFF1;
    // rom_array[19789] = 32'hFFFFFFF0;
    // rom_array[19790] = 32'hFFFFFFF0;
    // rom_array[19791] = 32'hFFFFFFF1;
    // rom_array[19792] = 32'hFFFFFFF1;
    // rom_array[19793] = 32'hFFFFFFF0;
    // rom_array[19794] = 32'hFFFFFFF0;
    // rom_array[19795] = 32'hFFFFFFF1;
    // rom_array[19796] = 32'hFFFFFFF1;
    // rom_array[19797] = 32'hFFFFFFF0;
    // rom_array[19798] = 32'hFFFFFFF0;
    // rom_array[19799] = 32'hFFFFFFF1;
    // rom_array[19800] = 32'hFFFFFFF1;
    // rom_array[19801] = 32'hFFFFFFF0;
    // rom_array[19802] = 32'hFFFFFFF0;
    // rom_array[19803] = 32'hFFFFFFF1;
    // rom_array[19804] = 32'hFFFFFFF1;
    // rom_array[19805] = 32'hFFFFFFF0;
    // rom_array[19806] = 32'hFFFFFFF0;
    // rom_array[19807] = 32'hFFFFFFF1;
    // rom_array[19808] = 32'hFFFFFFF1;
    // rom_array[19809] = 32'hFFFFFFF0;
    // rom_array[19810] = 32'hFFFFFFF0;
    // rom_array[19811] = 32'hFFFFFFF1;
    // rom_array[19812] = 32'hFFFFFFF1;
    // rom_array[19813] = 32'hFFFFFFF0;
    // rom_array[19814] = 32'hFFFFFFF0;
    // rom_array[19815] = 32'hFFFFFFF1;
    // rom_array[19816] = 32'hFFFFFFF1;
    // rom_array[19817] = 32'hFFFFFFF0;
    // rom_array[19818] = 32'hFFFFFFF0;
    // rom_array[19819] = 32'hFFFFFFF1;
    // rom_array[19820] = 32'hFFFFFFF1;
    // rom_array[19821] = 32'hFFFFFFF0;
    // rom_array[19822] = 32'hFFFFFFF0;
    // rom_array[19823] = 32'hFFFFFFF1;
    // rom_array[19824] = 32'hFFFFFFF1;
    // rom_array[19825] = 32'hFFFFFFF0;
    // rom_array[19826] = 32'hFFFFFFF0;
    // rom_array[19827] = 32'hFFFFFFF1;
    // rom_array[19828] = 32'hFFFFFFF1;
    // rom_array[19829] = 32'hFFFFFFF0;
    // rom_array[19830] = 32'hFFFFFFF0;
    // rom_array[19831] = 32'hFFFFFFF1;
    // rom_array[19832] = 32'hFFFFFFF1;
    // rom_array[19833] = 32'hFFFFFFF0;
    // rom_array[19834] = 32'hFFFFFFF0;
    // rom_array[19835] = 32'hFFFFFFF1;
    // rom_array[19836] = 32'hFFFFFFF1;
    // rom_array[19837] = 32'hFFFFFFF0;
    // rom_array[19838] = 32'hFFFFFFF0;
    // rom_array[19839] = 32'hFFFFFFF1;
    // rom_array[19840] = 32'hFFFFFFF1;
    // rom_array[19841] = 32'hFFFFFFF0;
    // rom_array[19842] = 32'hFFFFFFF0;
    // rom_array[19843] = 32'hFFFFFFF1;
    // rom_array[19844] = 32'hFFFFFFF1;
    // rom_array[19845] = 32'hFFFFFFF0;
    // rom_array[19846] = 32'hFFFFFFF0;
    // rom_array[19847] = 32'hFFFFFFF1;
    // rom_array[19848] = 32'hFFFFFFF1;
    // rom_array[19849] = 32'hFFFFFFF0;
    // rom_array[19850] = 32'hFFFFFFF0;
    // rom_array[19851] = 32'hFFFFFFF1;
    // rom_array[19852] = 32'hFFFFFFF1;
    // rom_array[19853] = 32'hFFFFFFF0;
    // rom_array[19854] = 32'hFFFFFFF0;
    // rom_array[19855] = 32'hFFFFFFF1;
    // rom_array[19856] = 32'hFFFFFFF1;
    // rom_array[19857] = 32'hFFFFFFF0;
    // rom_array[19858] = 32'hFFFFFFF0;
    // rom_array[19859] = 32'hFFFFFFF1;
    // rom_array[19860] = 32'hFFFFFFF1;
    // rom_array[19861] = 32'hFFFFFFF0;
    // rom_array[19862] = 32'hFFFFFFF0;
    // rom_array[19863] = 32'hFFFFFFF1;
    // rom_array[19864] = 32'hFFFFFFF1;
    // rom_array[19865] = 32'hFFFFFFF0;
    // rom_array[19866] = 32'hFFFFFFF0;
    // rom_array[19867] = 32'hFFFFFFF0;
    // rom_array[19868] = 32'hFFFFFFF0;
    // rom_array[19869] = 32'hFFFFFFF0;
    // rom_array[19870] = 32'hFFFFFFF0;
    // rom_array[19871] = 32'hFFFFFFF1;
    // rom_array[19872] = 32'hFFFFFFF1;
    // rom_array[19873] = 32'hFFFFFFF0;
    // rom_array[19874] = 32'hFFFFFFF0;
    // rom_array[19875] = 32'hFFFFFFF0;
    // rom_array[19876] = 32'hFFFFFFF0;
    // rom_array[19877] = 32'hFFFFFFF0;
    // rom_array[19878] = 32'hFFFFFFF0;
    // rom_array[19879] = 32'hFFFFFFF1;
    // rom_array[19880] = 32'hFFFFFFF1;
    // rom_array[19881] = 32'hFFFFFFF0;
    // rom_array[19882] = 32'hFFFFFFF0;
    // rom_array[19883] = 32'hFFFFFFF1;
    // rom_array[19884] = 32'hFFFFFFF1;
    // rom_array[19885] = 32'hFFFFFFF0;
    // rom_array[19886] = 32'hFFFFFFF0;
    // rom_array[19887] = 32'hFFFFFFF0;
    // rom_array[19888] = 32'hFFFFFFF0;
    // rom_array[19889] = 32'hFFFFFFF0;
    // rom_array[19890] = 32'hFFFFFFF0;
    // rom_array[19891] = 32'hFFFFFFF1;
    // rom_array[19892] = 32'hFFFFFFF1;
    // rom_array[19893] = 32'hFFFFFFF0;
    // rom_array[19894] = 32'hFFFFFFF0;
    // rom_array[19895] = 32'hFFFFFFF0;
    // rom_array[19896] = 32'hFFFFFFF0;
    // rom_array[19897] = 32'hFFFFFFF1;
    // rom_array[19898] = 32'hFFFFFFF1;
    // rom_array[19899] = 32'hFFFFFFF1;
    // rom_array[19900] = 32'hFFFFFFF1;
    // rom_array[19901] = 32'hFFFFFFF0;
    // rom_array[19902] = 32'hFFFFFFF0;
    // rom_array[19903] = 32'hFFFFFFF0;
    // rom_array[19904] = 32'hFFFFFFF0;
    // rom_array[19905] = 32'hFFFFFFF1;
    // rom_array[19906] = 32'hFFFFFFF1;
    // rom_array[19907] = 32'hFFFFFFF1;
    // rom_array[19908] = 32'hFFFFFFF1;
    // rom_array[19909] = 32'hFFFFFFF0;
    // rom_array[19910] = 32'hFFFFFFF0;
    // rom_array[19911] = 32'hFFFFFFF0;
    // rom_array[19912] = 32'hFFFFFFF0;
    // rom_array[19913] = 32'hFFFFFFF1;
    // rom_array[19914] = 32'hFFFFFFF1;
    // rom_array[19915] = 32'hFFFFFFF1;
    // rom_array[19916] = 32'hFFFFFFF1;
    // rom_array[19917] = 32'hFFFFFFF0;
    // rom_array[19918] = 32'hFFFFFFF0;
    // rom_array[19919] = 32'hFFFFFFF0;
    // rom_array[19920] = 32'hFFFFFFF0;
    // rom_array[19921] = 32'hFFFFFFF1;
    // rom_array[19922] = 32'hFFFFFFF1;
    // rom_array[19923] = 32'hFFFFFFF1;
    // rom_array[19924] = 32'hFFFFFFF1;
    // rom_array[19925] = 32'hFFFFFFF0;
    // rom_array[19926] = 32'hFFFFFFF0;
    // rom_array[19927] = 32'hFFFFFFF0;
    // rom_array[19928] = 32'hFFFFFFF0;
    // rom_array[19929] = 32'hFFFFFFF1;
    // rom_array[19930] = 32'hFFFFFFF1;
    // rom_array[19931] = 32'hFFFFFFF1;
    // rom_array[19932] = 32'hFFFFFFF1;
    // rom_array[19933] = 32'hFFFFFFF0;
    // rom_array[19934] = 32'hFFFFFFF0;
    // rom_array[19935] = 32'hFFFFFFF1;
    // rom_array[19936] = 32'hFFFFFFF1;
    // rom_array[19937] = 32'hFFFFFFF1;
    // rom_array[19938] = 32'hFFFFFFF1;
    // rom_array[19939] = 32'hFFFFFFF1;
    // rom_array[19940] = 32'hFFFFFFF1;
    // rom_array[19941] = 32'hFFFFFFF0;
    // rom_array[19942] = 32'hFFFFFFF0;
    // rom_array[19943] = 32'hFFFFFFF1;
    // rom_array[19944] = 32'hFFFFFFF1;
    // rom_array[19945] = 32'hFFFFFFF0;
    // rom_array[19946] = 32'hFFFFFFF0;
    // rom_array[19947] = 32'hFFFFFFF1;
    // rom_array[19948] = 32'hFFFFFFF1;
    // rom_array[19949] = 32'hFFFFFFF0;
    // rom_array[19950] = 32'hFFFFFFF0;
    // rom_array[19951] = 32'hFFFFFFF1;
    // rom_array[19952] = 32'hFFFFFFF1;
    // rom_array[19953] = 32'hFFFFFFF0;
    // rom_array[19954] = 32'hFFFFFFF0;
    // rom_array[19955] = 32'hFFFFFFF1;
    // rom_array[19956] = 32'hFFFFFFF1;
    // rom_array[19957] = 32'hFFFFFFF0;
    // rom_array[19958] = 32'hFFFFFFF0;
    // rom_array[19959] = 32'hFFFFFFF1;
    // rom_array[19960] = 32'hFFFFFFF1;
    // rom_array[19961] = 32'hFFFFFFF0;
    // rom_array[19962] = 32'hFFFFFFF0;
    // rom_array[19963] = 32'hFFFFFFF1;
    // rom_array[19964] = 32'hFFFFFFF1;
    // rom_array[19965] = 32'hFFFFFFF0;
    // rom_array[19966] = 32'hFFFFFFF0;
    // rom_array[19967] = 32'hFFFFFFF1;
    // rom_array[19968] = 32'hFFFFFFF1;
    // rom_array[19969] = 32'hFFFFFFF0;
    // rom_array[19970] = 32'hFFFFFFF0;
    // rom_array[19971] = 32'hFFFFFFF1;
    // rom_array[19972] = 32'hFFFFFFF1;
    // rom_array[19973] = 32'hFFFFFFF0;
    // rom_array[19974] = 32'hFFFFFFF0;
    // rom_array[19975] = 32'hFFFFFFF1;
    // rom_array[19976] = 32'hFFFFFFF1;
    // rom_array[19977] = 32'hFFFFFFF0;
    // rom_array[19978] = 32'hFFFFFFF0;
    // rom_array[19979] = 32'hFFFFFFF1;
    // rom_array[19980] = 32'hFFFFFFF1;
    // rom_array[19981] = 32'hFFFFFFF0;
    // rom_array[19982] = 32'hFFFFFFF0;
    // rom_array[19983] = 32'hFFFFFFF0;
    // rom_array[19984] = 32'hFFFFFFF0;
    // rom_array[19985] = 32'hFFFFFFF0;
    // rom_array[19986] = 32'hFFFFFFF0;
    // rom_array[19987] = 32'hFFFFFFF1;
    // rom_array[19988] = 32'hFFFFFFF1;
    // rom_array[19989] = 32'hFFFFFFF0;
    // rom_array[19990] = 32'hFFFFFFF0;
    // rom_array[19991] = 32'hFFFFFFF0;
    // rom_array[19992] = 32'hFFFFFFF0;
    // rom_array[19993] = 32'hFFFFFFF0;
    // rom_array[19994] = 32'hFFFFFFF0;
    // rom_array[19995] = 32'hFFFFFFF0;
    // rom_array[19996] = 32'hFFFFFFF0;
    // rom_array[19997] = 32'hFFFFFFF0;
    // rom_array[19998] = 32'hFFFFFFF0;
    // rom_array[19999] = 32'hFFFFFFF1;
    // rom_array[20000] = 32'hFFFFFFF1;
    // rom_array[20001] = 32'hFFFFFFF0;
    // rom_array[20002] = 32'hFFFFFFF0;
    // rom_array[20003] = 32'hFFFFFFF0;
    // rom_array[20004] = 32'hFFFFFFF0;
    // rom_array[20005] = 32'hFFFFFFF0;
    // rom_array[20006] = 32'hFFFFFFF0;
    // rom_array[20007] = 32'hFFFFFFF1;
    // rom_array[20008] = 32'hFFFFFFF1;
    // rom_array[20009] = 32'hFFFFFFF0;
    // rom_array[20010] = 32'hFFFFFFF0;
    // rom_array[20011] = 32'hFFFFFFF0;
    // rom_array[20012] = 32'hFFFFFFF0;
    // rom_array[20013] = 32'hFFFFFFF1;
    // rom_array[20014] = 32'hFFFFFFF1;
    // rom_array[20015] = 32'hFFFFFFF1;
    // rom_array[20016] = 32'hFFFFFFF1;
    // rom_array[20017] = 32'hFFFFFFF0;
    // rom_array[20018] = 32'hFFFFFFF0;
    // rom_array[20019] = 32'hFFFFFFF0;
    // rom_array[20020] = 32'hFFFFFFF0;
    // rom_array[20021] = 32'hFFFFFFF1;
    // rom_array[20022] = 32'hFFFFFFF1;
    // rom_array[20023] = 32'hFFFFFFF1;
    // rom_array[20024] = 32'hFFFFFFF1;
    // rom_array[20025] = 32'hFFFFFFF0;
    // rom_array[20026] = 32'hFFFFFFF0;
    // rom_array[20027] = 32'hFFFFFFF1;
    // rom_array[20028] = 32'hFFFFFFF1;
    // rom_array[20029] = 32'hFFFFFFF0;
    // rom_array[20030] = 32'hFFFFFFF0;
    // rom_array[20031] = 32'hFFFFFFF1;
    // rom_array[20032] = 32'hFFFFFFF1;
    // rom_array[20033] = 32'hFFFFFFF0;
    // rom_array[20034] = 32'hFFFFFFF0;
    // rom_array[20035] = 32'hFFFFFFF1;
    // rom_array[20036] = 32'hFFFFFFF1;
    // rom_array[20037] = 32'hFFFFFFF0;
    // rom_array[20038] = 32'hFFFFFFF0;
    // rom_array[20039] = 32'hFFFFFFF1;
    // rom_array[20040] = 32'hFFFFFFF1;
    // rom_array[20041] = 32'hFFFFFFF0;
    // rom_array[20042] = 32'hFFFFFFF0;
    // rom_array[20043] = 32'hFFFFFFF0;
    // rom_array[20044] = 32'hFFFFFFF0;
    // rom_array[20045] = 32'hFFFFFFF1;
    // rom_array[20046] = 32'hFFFFFFF1;
    // rom_array[20047] = 32'hFFFFFFF1;
    // rom_array[20048] = 32'hFFFFFFF1;
    // rom_array[20049] = 32'hFFFFFFF0;
    // rom_array[20050] = 32'hFFFFFFF0;
    // rom_array[20051] = 32'hFFFFFFF0;
    // rom_array[20052] = 32'hFFFFFFF0;
    // rom_array[20053] = 32'hFFFFFFF1;
    // rom_array[20054] = 32'hFFFFFFF1;
    // rom_array[20055] = 32'hFFFFFFF1;
    // rom_array[20056] = 32'hFFFFFFF1;
    // rom_array[20057] = 32'hFFFFFFF0;
    // rom_array[20058] = 32'hFFFFFFF0;
    // rom_array[20059] = 32'hFFFFFFF0;
    // rom_array[20060] = 32'hFFFFFFF0;
    // rom_array[20061] = 32'hFFFFFFF1;
    // rom_array[20062] = 32'hFFFFFFF1;
    // rom_array[20063] = 32'hFFFFFFF1;
    // rom_array[20064] = 32'hFFFFFFF1;
    // rom_array[20065] = 32'hFFFFFFF0;
    // rom_array[20066] = 32'hFFFFFFF0;
    // rom_array[20067] = 32'hFFFFFFF0;
    // rom_array[20068] = 32'hFFFFFFF0;
    // rom_array[20069] = 32'hFFFFFFF1;
    // rom_array[20070] = 32'hFFFFFFF1;
    // rom_array[20071] = 32'hFFFFFFF1;
    // rom_array[20072] = 32'hFFFFFFF1;
    // rom_array[20073] = 32'hFFFFFFF0;
    // rom_array[20074] = 32'hFFFFFFF0;
    // rom_array[20075] = 32'hFFFFFFF1;
    // rom_array[20076] = 32'hFFFFFFF1;
    // rom_array[20077] = 32'hFFFFFFF0;
    // rom_array[20078] = 32'hFFFFFFF0;
    // rom_array[20079] = 32'hFFFFFFF1;
    // rom_array[20080] = 32'hFFFFFFF1;
    // rom_array[20081] = 32'hFFFFFFF0;
    // rom_array[20082] = 32'hFFFFFFF0;
    // rom_array[20083] = 32'hFFFFFFF1;
    // rom_array[20084] = 32'hFFFFFFF1;
    // rom_array[20085] = 32'hFFFFFFF0;
    // rom_array[20086] = 32'hFFFFFFF0;
    // rom_array[20087] = 32'hFFFFFFF1;
    // rom_array[20088] = 32'hFFFFFFF1;
    // rom_array[20089] = 32'hFFFFFFF0;
    // rom_array[20090] = 32'hFFFFFFF0;
    // rom_array[20091] = 32'hFFFFFFF1;
    // rom_array[20092] = 32'hFFFFFFF1;
    // rom_array[20093] = 32'hFFFFFFF0;
    // rom_array[20094] = 32'hFFFFFFF0;
    // rom_array[20095] = 32'hFFFFFFF1;
    // rom_array[20096] = 32'hFFFFFFF1;
    // rom_array[20097] = 32'hFFFFFFF0;
    // rom_array[20098] = 32'hFFFFFFF0;
    // rom_array[20099] = 32'hFFFFFFF1;
    // rom_array[20100] = 32'hFFFFFFF1;
    // rom_array[20101] = 32'hFFFFFFF0;
    // rom_array[20102] = 32'hFFFFFFF0;
    // rom_array[20103] = 32'hFFFFFFF1;
    // rom_array[20104] = 32'hFFFFFFF1;
    // rom_array[20105] = 32'hFFFFFFF0;
    // rom_array[20106] = 32'hFFFFFFF0;
    // rom_array[20107] = 32'hFFFFFFF1;
    // rom_array[20108] = 32'hFFFFFFF1;
    // rom_array[20109] = 32'hFFFFFFF0;
    // rom_array[20110] = 32'hFFFFFFF0;
    // rom_array[20111] = 32'hFFFFFFF1;
    // rom_array[20112] = 32'hFFFFFFF1;
    // rom_array[20113] = 32'hFFFFFFF0;
    // rom_array[20114] = 32'hFFFFFFF0;
    // rom_array[20115] = 32'hFFFFFFF1;
    // rom_array[20116] = 32'hFFFFFFF1;
    // rom_array[20117] = 32'hFFFFFFF0;
    // rom_array[20118] = 32'hFFFFFFF0;
    // rom_array[20119] = 32'hFFFFFFF1;
    // rom_array[20120] = 32'hFFFFFFF1;
    // rom_array[20121] = 32'hFFFFFFF1;
    // rom_array[20122] = 32'hFFFFFFF1;
    // rom_array[20123] = 32'hFFFFFFF1;
    // rom_array[20124] = 32'hFFFFFFF1;
    // rom_array[20125] = 32'hFFFFFFF1;
    // rom_array[20126] = 32'hFFFFFFF1;
    // rom_array[20127] = 32'hFFFFFFF1;
    // rom_array[20128] = 32'hFFFFFFF1;
    // rom_array[20129] = 32'hFFFFFFF1;
    // rom_array[20130] = 32'hFFFFFFF1;
    // rom_array[20131] = 32'hFFFFFFF1;
    // rom_array[20132] = 32'hFFFFFFF1;
    // rom_array[20133] = 32'hFFFFFFF1;
    // rom_array[20134] = 32'hFFFFFFF1;
    // rom_array[20135] = 32'hFFFFFFF1;
    // rom_array[20136] = 32'hFFFFFFF1;
    // rom_array[20137] = 32'hFFFFFFF0;
    // rom_array[20138] = 32'hFFFFFFF0;
    // rom_array[20139] = 32'hFFFFFFF1;
    // rom_array[20140] = 32'hFFFFFFF1;
    // rom_array[20141] = 32'hFFFFFFF0;
    // rom_array[20142] = 32'hFFFFFFF0;
    // rom_array[20143] = 32'hFFFFFFF1;
    // rom_array[20144] = 32'hFFFFFFF1;
    // rom_array[20145] = 32'hFFFFFFF0;
    // rom_array[20146] = 32'hFFFFFFF0;
    // rom_array[20147] = 32'hFFFFFFF1;
    // rom_array[20148] = 32'hFFFFFFF1;
    // rom_array[20149] = 32'hFFFFFFF0;
    // rom_array[20150] = 32'hFFFFFFF0;
    // rom_array[20151] = 32'hFFFFFFF1;
    // rom_array[20152] = 32'hFFFFFFF1;
    // rom_array[20153] = 32'hFFFFFFF1;
    // rom_array[20154] = 32'hFFFFFFF1;
    // rom_array[20155] = 32'hFFFFFFF1;
    // rom_array[20156] = 32'hFFFFFFF1;
    // rom_array[20157] = 32'hFFFFFFF1;
    // rom_array[20158] = 32'hFFFFFFF1;
    // rom_array[20159] = 32'hFFFFFFF1;
    // rom_array[20160] = 32'hFFFFFFF1;
    // rom_array[20161] = 32'hFFFFFFF1;
    // rom_array[20162] = 32'hFFFFFFF1;
    // rom_array[20163] = 32'hFFFFFFF1;
    // rom_array[20164] = 32'hFFFFFFF1;
    // rom_array[20165] = 32'hFFFFFFF1;
    // rom_array[20166] = 32'hFFFFFFF1;
    // rom_array[20167] = 32'hFFFFFFF1;
    // rom_array[20168] = 32'hFFFFFFF1;
    // rom_array[20169] = 32'hFFFFFFF1;
    // rom_array[20170] = 32'hFFFFFFF1;
    // rom_array[20171] = 32'hFFFFFFF1;
    // rom_array[20172] = 32'hFFFFFFF1;
    // rom_array[20173] = 32'hFFFFFFF1;
    // rom_array[20174] = 32'hFFFFFFF1;
    // rom_array[20175] = 32'hFFFFFFF1;
    // rom_array[20176] = 32'hFFFFFFF1;
    // rom_array[20177] = 32'hFFFFFFF1;
    // rom_array[20178] = 32'hFFFFFFF1;
    // rom_array[20179] = 32'hFFFFFFF1;
    // rom_array[20180] = 32'hFFFFFFF1;
    // rom_array[20181] = 32'hFFFFFFF1;
    // rom_array[20182] = 32'hFFFFFFF1;
    // rom_array[20183] = 32'hFFFFFFF1;
    // rom_array[20184] = 32'hFFFFFFF1;
    // rom_array[20185] = 32'hFFFFFFF0;
    // rom_array[20186] = 32'hFFFFFFF0;
    // rom_array[20187] = 32'hFFFFFFF0;
    // rom_array[20188] = 32'hFFFFFFF0;
    // rom_array[20189] = 32'hFFFFFFF1;
    // rom_array[20190] = 32'hFFFFFFF1;
    // rom_array[20191] = 32'hFFFFFFF1;
    // rom_array[20192] = 32'hFFFFFFF1;
    // rom_array[20193] = 32'hFFFFFFF0;
    // rom_array[20194] = 32'hFFFFFFF0;
    // rom_array[20195] = 32'hFFFFFFF0;
    // rom_array[20196] = 32'hFFFFFFF0;
    // rom_array[20197] = 32'hFFFFFFF1;
    // rom_array[20198] = 32'hFFFFFFF1;
    // rom_array[20199] = 32'hFFFFFFF1;
    // rom_array[20200] = 32'hFFFFFFF1;
    // rom_array[20201] = 32'hFFFFFFF0;
    // rom_array[20202] = 32'hFFFFFFF0;
    // rom_array[20203] = 32'hFFFFFFF0;
    // rom_array[20204] = 32'hFFFFFFF0;
    // rom_array[20205] = 32'hFFFFFFF1;
    // rom_array[20206] = 32'hFFFFFFF1;
    // rom_array[20207] = 32'hFFFFFFF1;
    // rom_array[20208] = 32'hFFFFFFF1;
    // rom_array[20209] = 32'hFFFFFFF0;
    // rom_array[20210] = 32'hFFFFFFF0;
    // rom_array[20211] = 32'hFFFFFFF0;
    // rom_array[20212] = 32'hFFFFFFF0;
    // rom_array[20213] = 32'hFFFFFFF1;
    // rom_array[20214] = 32'hFFFFFFF1;
    // rom_array[20215] = 32'hFFFFFFF1;
    // rom_array[20216] = 32'hFFFFFFF1;
    // rom_array[20217] = 32'hFFFFFFF0;
    // rom_array[20218] = 32'hFFFFFFF0;
    // rom_array[20219] = 32'hFFFFFFF0;
    // rom_array[20220] = 32'hFFFFFFF0;
    // rom_array[20221] = 32'hFFFFFFF1;
    // rom_array[20222] = 32'hFFFFFFF1;
    // rom_array[20223] = 32'hFFFFFFF1;
    // rom_array[20224] = 32'hFFFFFFF1;
    // rom_array[20225] = 32'hFFFFFFF0;
    // rom_array[20226] = 32'hFFFFFFF0;
    // rom_array[20227] = 32'hFFFFFFF0;
    // rom_array[20228] = 32'hFFFFFFF0;
    // rom_array[20229] = 32'hFFFFFFF1;
    // rom_array[20230] = 32'hFFFFFFF1;
    // rom_array[20231] = 32'hFFFFFFF1;
    // rom_array[20232] = 32'hFFFFFFF1;
    // rom_array[20233] = 32'hFFFFFFF0;
    // rom_array[20234] = 32'hFFFFFFF0;
    // rom_array[20235] = 32'hFFFFFFF0;
    // rom_array[20236] = 32'hFFFFFFF0;
    // rom_array[20237] = 32'hFFFFFFF1;
    // rom_array[20238] = 32'hFFFFFFF1;
    // rom_array[20239] = 32'hFFFFFFF1;
    // rom_array[20240] = 32'hFFFFFFF1;
    // rom_array[20241] = 32'hFFFFFFF0;
    // rom_array[20242] = 32'hFFFFFFF0;
    // rom_array[20243] = 32'hFFFFFFF0;
    // rom_array[20244] = 32'hFFFFFFF0;
    // rom_array[20245] = 32'hFFFFFFF1;
    // rom_array[20246] = 32'hFFFFFFF1;
    // rom_array[20247] = 32'hFFFFFFF1;
    // rom_array[20248] = 32'hFFFFFFF1;
    // rom_array[20249] = 32'hFFFFFFF0;
    // rom_array[20250] = 32'hFFFFFFF0;
    // rom_array[20251] = 32'hFFFFFFF0;
    // rom_array[20252] = 32'hFFFFFFF0;
    // rom_array[20253] = 32'hFFFFFFF1;
    // rom_array[20254] = 32'hFFFFFFF1;
    // rom_array[20255] = 32'hFFFFFFF1;
    // rom_array[20256] = 32'hFFFFFFF1;
    // rom_array[20257] = 32'hFFFFFFF0;
    // rom_array[20258] = 32'hFFFFFFF0;
    // rom_array[20259] = 32'hFFFFFFF0;
    // rom_array[20260] = 32'hFFFFFFF0;
    // rom_array[20261] = 32'hFFFFFFF1;
    // rom_array[20262] = 32'hFFFFFFF1;
    // rom_array[20263] = 32'hFFFFFFF1;
    // rom_array[20264] = 32'hFFFFFFF1;
    // rom_array[20265] = 32'hFFFFFFF0;
    // rom_array[20266] = 32'hFFFFFFF0;
    // rom_array[20267] = 32'hFFFFFFF0;
    // rom_array[20268] = 32'hFFFFFFF0;
    // rom_array[20269] = 32'hFFFFFFF1;
    // rom_array[20270] = 32'hFFFFFFF1;
    // rom_array[20271] = 32'hFFFFFFF1;
    // rom_array[20272] = 32'hFFFFFFF1;
    // rom_array[20273] = 32'hFFFFFFF0;
    // rom_array[20274] = 32'hFFFFFFF0;
    // rom_array[20275] = 32'hFFFFFFF0;
    // rom_array[20276] = 32'hFFFFFFF0;
    // rom_array[20277] = 32'hFFFFFFF1;
    // rom_array[20278] = 32'hFFFFFFF1;
    // rom_array[20279] = 32'hFFFFFFF1;
    // rom_array[20280] = 32'hFFFFFFF1;
    // rom_array[20281] = 32'hFFFFFFF0;
    // rom_array[20282] = 32'hFFFFFFF0;
    // rom_array[20283] = 32'hFFFFFFF0;
    // rom_array[20284] = 32'hFFFFFFF0;
    // rom_array[20285] = 32'hFFFFFFF1;
    // rom_array[20286] = 32'hFFFFFFF1;
    // rom_array[20287] = 32'hFFFFFFF1;
    // rom_array[20288] = 32'hFFFFFFF1;
    // rom_array[20289] = 32'hFFFFFFF0;
    // rom_array[20290] = 32'hFFFFFFF0;
    // rom_array[20291] = 32'hFFFFFFF0;
    // rom_array[20292] = 32'hFFFFFFF0;
    // rom_array[20293] = 32'hFFFFFFF1;
    // rom_array[20294] = 32'hFFFFFFF1;
    // rom_array[20295] = 32'hFFFFFFF1;
    // rom_array[20296] = 32'hFFFFFFF1;
    // rom_array[20297] = 32'hFFFFFFF0;
    // rom_array[20298] = 32'hFFFFFFF0;
    // rom_array[20299] = 32'hFFFFFFF0;
    // rom_array[20300] = 32'hFFFFFFF0;
    // rom_array[20301] = 32'hFFFFFFF1;
    // rom_array[20302] = 32'hFFFFFFF1;
    // rom_array[20303] = 32'hFFFFFFF1;
    // rom_array[20304] = 32'hFFFFFFF1;
    // rom_array[20305] = 32'hFFFFFFF0;
    // rom_array[20306] = 32'hFFFFFFF0;
    // rom_array[20307] = 32'hFFFFFFF0;
    // rom_array[20308] = 32'hFFFFFFF0;
    // rom_array[20309] = 32'hFFFFFFF1;
    // rom_array[20310] = 32'hFFFFFFF1;
    // rom_array[20311] = 32'hFFFFFFF1;
    // rom_array[20312] = 32'hFFFFFFF1;
    // rom_array[20313] = 32'hFFFFFFF1;
    // rom_array[20314] = 32'hFFFFFFF1;
    // rom_array[20315] = 32'hFFFFFFF1;
    // rom_array[20316] = 32'hFFFFFFF1;
    // rom_array[20317] = 32'hFFFFFFF1;
    // rom_array[20318] = 32'hFFFFFFF1;
    // rom_array[20319] = 32'hFFFFFFF1;
    // rom_array[20320] = 32'hFFFFFFF1;
    // rom_array[20321] = 32'hFFFFFFF1;
    // rom_array[20322] = 32'hFFFFFFF1;
    // rom_array[20323] = 32'hFFFFFFF1;
    // rom_array[20324] = 32'hFFFFFFF1;
    // rom_array[20325] = 32'hFFFFFFF1;
    // rom_array[20326] = 32'hFFFFFFF1;
    // rom_array[20327] = 32'hFFFFFFF1;
    // rom_array[20328] = 32'hFFFFFFF1;
    // rom_array[20329] = 32'hFFFFFFF1;
    // rom_array[20330] = 32'hFFFFFFF1;
    // rom_array[20331] = 32'hFFFFFFF1;
    // rom_array[20332] = 32'hFFFFFFF1;
    // rom_array[20333] = 32'hFFFFFFF0;
    // rom_array[20334] = 32'hFFFFFFF0;
    // rom_array[20335] = 32'hFFFFFFF0;
    // rom_array[20336] = 32'hFFFFFFF0;
    // rom_array[20337] = 32'hFFFFFFF1;
    // rom_array[20338] = 32'hFFFFFFF1;
    // rom_array[20339] = 32'hFFFFFFF1;
    // rom_array[20340] = 32'hFFFFFFF1;
    // rom_array[20341] = 32'hFFFFFFF0;
    // rom_array[20342] = 32'hFFFFFFF0;
    // rom_array[20343] = 32'hFFFFFFF0;
    // rom_array[20344] = 32'hFFFFFFF0;
    // rom_array[20345] = 32'hFFFFFFF1;
    // rom_array[20346] = 32'hFFFFFFF1;
    // rom_array[20347] = 32'hFFFFFFF1;
    // rom_array[20348] = 32'hFFFFFFF1;
    // rom_array[20349] = 32'hFFFFFFF1;
    // rom_array[20350] = 32'hFFFFFFF1;
    // rom_array[20351] = 32'hFFFFFFF1;
    // rom_array[20352] = 32'hFFFFFFF1;
    // rom_array[20353] = 32'hFFFFFFF1;
    // rom_array[20354] = 32'hFFFFFFF1;
    // rom_array[20355] = 32'hFFFFFFF1;
    // rom_array[20356] = 32'hFFFFFFF1;
    // rom_array[20357] = 32'hFFFFFFF1;
    // rom_array[20358] = 32'hFFFFFFF1;
    // rom_array[20359] = 32'hFFFFFFF1;
    // rom_array[20360] = 32'hFFFFFFF1;
    // rom_array[20361] = 32'hFFFFFFF1;
    // rom_array[20362] = 32'hFFFFFFF1;
    // rom_array[20363] = 32'hFFFFFFF1;
    // rom_array[20364] = 32'hFFFFFFF1;
    // rom_array[20365] = 32'hFFFFFFF0;
    // rom_array[20366] = 32'hFFFFFFF0;
    // rom_array[20367] = 32'hFFFFFFF0;
    // rom_array[20368] = 32'hFFFFFFF0;
    // rom_array[20369] = 32'hFFFFFFF1;
    // rom_array[20370] = 32'hFFFFFFF1;
    // rom_array[20371] = 32'hFFFFFFF1;
    // rom_array[20372] = 32'hFFFFFFF1;
    // rom_array[20373] = 32'hFFFFFFF0;
    // rom_array[20374] = 32'hFFFFFFF0;
    // rom_array[20375] = 32'hFFFFFFF0;
    // rom_array[20376] = 32'hFFFFFFF0;
    // rom_array[20377] = 32'hFFFFFFF1;
    // rom_array[20378] = 32'hFFFFFFF1;
    // rom_array[20379] = 32'hFFFFFFF1;
    // rom_array[20380] = 32'hFFFFFFF1;
    // rom_array[20381] = 32'hFFFFFFF0;
    // rom_array[20382] = 32'hFFFFFFF0;
    // rom_array[20383] = 32'hFFFFFFF0;
    // rom_array[20384] = 32'hFFFFFFF0;
    // rom_array[20385] = 32'hFFFFFFF1;
    // rom_array[20386] = 32'hFFFFFFF1;
    // rom_array[20387] = 32'hFFFFFFF1;
    // rom_array[20388] = 32'hFFFFFFF1;
    // rom_array[20389] = 32'hFFFFFFF0;
    // rom_array[20390] = 32'hFFFFFFF0;
    // rom_array[20391] = 32'hFFFFFFF0;
    // rom_array[20392] = 32'hFFFFFFF0;
    // rom_array[20393] = 32'hFFFFFFF1;
    // rom_array[20394] = 32'hFFFFFFF1;
    // rom_array[20395] = 32'hFFFFFFF1;
    // rom_array[20396] = 32'hFFFFFFF1;
    // rom_array[20397] = 32'hFFFFFFF0;
    // rom_array[20398] = 32'hFFFFFFF0;
    // rom_array[20399] = 32'hFFFFFFF0;
    // rom_array[20400] = 32'hFFFFFFF0;
    // rom_array[20401] = 32'hFFFFFFF1;
    // rom_array[20402] = 32'hFFFFFFF1;
    // rom_array[20403] = 32'hFFFFFFF1;
    // rom_array[20404] = 32'hFFFFFFF1;
    // rom_array[20405] = 32'hFFFFFFF0;
    // rom_array[20406] = 32'hFFFFFFF0;
    // rom_array[20407] = 32'hFFFFFFF0;
    // rom_array[20408] = 32'hFFFFFFF0;
    // rom_array[20409] = 32'hFFFFFFF1;
    // rom_array[20410] = 32'hFFFFFFF1;
    // rom_array[20411] = 32'hFFFFFFF1;
    // rom_array[20412] = 32'hFFFFFFF1;
    // rom_array[20413] = 32'hFFFFFFF0;
    // rom_array[20414] = 32'hFFFFFFF0;
    // rom_array[20415] = 32'hFFFFFFF1;
    // rom_array[20416] = 32'hFFFFFFF1;
    // rom_array[20417] = 32'hFFFFFFF1;
    // rom_array[20418] = 32'hFFFFFFF1;
    // rom_array[20419] = 32'hFFFFFFF1;
    // rom_array[20420] = 32'hFFFFFFF1;
    // rom_array[20421] = 32'hFFFFFFF0;
    // rom_array[20422] = 32'hFFFFFFF0;
    // rom_array[20423] = 32'hFFFFFFF1;
    // rom_array[20424] = 32'hFFFFFFF1;
    // rom_array[20425] = 32'hFFFFFFF0;
    // rom_array[20426] = 32'hFFFFFFF0;
    // rom_array[20427] = 32'hFFFFFFF1;
    // rom_array[20428] = 32'hFFFFFFF1;
    // rom_array[20429] = 32'hFFFFFFF0;
    // rom_array[20430] = 32'hFFFFFFF0;
    // rom_array[20431] = 32'hFFFFFFF1;
    // rom_array[20432] = 32'hFFFFFFF1;
    // rom_array[20433] = 32'hFFFFFFF0;
    // rom_array[20434] = 32'hFFFFFFF0;
    // rom_array[20435] = 32'hFFFFFFF1;
    // rom_array[20436] = 32'hFFFFFFF1;
    // rom_array[20437] = 32'hFFFFFFF0;
    // rom_array[20438] = 32'hFFFFFFF0;
    // rom_array[20439] = 32'hFFFFFFF1;
    // rom_array[20440] = 32'hFFFFFFF1;
    // rom_array[20441] = 32'hFFFFFFF1;
    // rom_array[20442] = 32'hFFFFFFF1;
    // rom_array[20443] = 32'hFFFFFFF1;
    // rom_array[20444] = 32'hFFFFFFF1;
    // rom_array[20445] = 32'hFFFFFFF1;
    // rom_array[20446] = 32'hFFFFFFF1;
    // rom_array[20447] = 32'hFFFFFFF1;
    // rom_array[20448] = 32'hFFFFFFF1;
    // rom_array[20449] = 32'hFFFFFFF1;
    // rom_array[20450] = 32'hFFFFFFF1;
    // rom_array[20451] = 32'hFFFFFFF1;
    // rom_array[20452] = 32'hFFFFFFF1;
    // rom_array[20453] = 32'hFFFFFFF1;
    // rom_array[20454] = 32'hFFFFFFF1;
    // rom_array[20455] = 32'hFFFFFFF1;
    // rom_array[20456] = 32'hFFFFFFF1;
    // rom_array[20457] = 32'hFFFFFFF1;
    // rom_array[20458] = 32'hFFFFFFF1;
    // rom_array[20459] = 32'hFFFFFFF1;
    // rom_array[20460] = 32'hFFFFFFF1;
    // rom_array[20461] = 32'hFFFFFFF1;
    // rom_array[20462] = 32'hFFFFFFF1;
    // rom_array[20463] = 32'hFFFFFFF1;
    // rom_array[20464] = 32'hFFFFFFF1;
    // rom_array[20465] = 32'hFFFFFFF1;
    // rom_array[20466] = 32'hFFFFFFF1;
    // rom_array[20467] = 32'hFFFFFFF1;
    // rom_array[20468] = 32'hFFFFFFF1;
    // rom_array[20469] = 32'hFFFFFFF1;
    // rom_array[20470] = 32'hFFFFFFF1;
    // rom_array[20471] = 32'hFFFFFFF1;
    // rom_array[20472] = 32'hFFFFFFF1;
    // rom_array[20473] = 32'hFFFFFFF0;
    // rom_array[20474] = 32'hFFFFFFF0;
    // rom_array[20475] = 32'hFFFFFFF1;
    // rom_array[20476] = 32'hFFFFFFF1;
    // rom_array[20477] = 32'hFFFFFFF0;
    // rom_array[20478] = 32'hFFFFFFF0;
    // rom_array[20479] = 32'hFFFFFFF1;
    // rom_array[20480] = 32'hFFFFFFF1;
    // rom_array[20481] = 32'hFFFFFFF0;
    // rom_array[20482] = 32'hFFFFFFF0;
    // rom_array[20483] = 32'hFFFFFFF1;
    // rom_array[20484] = 32'hFFFFFFF1;
    // rom_array[20485] = 32'hFFFFFFF0;
    // rom_array[20486] = 32'hFFFFFFF0;
    // rom_array[20487] = 32'hFFFFFFF1;
    // rom_array[20488] = 32'hFFFFFFF1;
    // rom_array[20489] = 32'hFFFFFFF0;
    // rom_array[20490] = 32'hFFFFFFF0;
    // rom_array[20491] = 32'hFFFFFFF1;
    // rom_array[20492] = 32'hFFFFFFF1;
    // rom_array[20493] = 32'hFFFFFFF0;
    // rom_array[20494] = 32'hFFFFFFF0;
    // rom_array[20495] = 32'hFFFFFFF1;
    // rom_array[20496] = 32'hFFFFFFF1;
    // rom_array[20497] = 32'hFFFFFFF0;
    // rom_array[20498] = 32'hFFFFFFF0;
    // rom_array[20499] = 32'hFFFFFFF1;
    // rom_array[20500] = 32'hFFFFFFF1;
    // rom_array[20501] = 32'hFFFFFFF0;
    // rom_array[20502] = 32'hFFFFFFF0;
    // rom_array[20503] = 32'hFFFFFFF1;
    // rom_array[20504] = 32'hFFFFFFF1;
    // rom_array[20505] = 32'hFFFFFFF0;
    // rom_array[20506] = 32'hFFFFFFF0;
    // rom_array[20507] = 32'hFFFFFFF1;
    // rom_array[20508] = 32'hFFFFFFF1;
    // rom_array[20509] = 32'hFFFFFFF0;
    // rom_array[20510] = 32'hFFFFFFF0;
    // rom_array[20511] = 32'hFFFFFFF1;
    // rom_array[20512] = 32'hFFFFFFF1;
    // rom_array[20513] = 32'hFFFFFFF0;
    // rom_array[20514] = 32'hFFFFFFF0;
    // rom_array[20515] = 32'hFFFFFFF1;
    // rom_array[20516] = 32'hFFFFFFF1;
    // rom_array[20517] = 32'hFFFFFFF0;
    // rom_array[20518] = 32'hFFFFFFF0;
    // rom_array[20519] = 32'hFFFFFFF1;
    // rom_array[20520] = 32'hFFFFFFF1;
    // rom_array[20521] = 32'hFFFFFFF0;
    // rom_array[20522] = 32'hFFFFFFF0;
    // rom_array[20523] = 32'hFFFFFFF1;
    // rom_array[20524] = 32'hFFFFFFF1;
    // rom_array[20525] = 32'hFFFFFFF0;
    // rom_array[20526] = 32'hFFFFFFF0;
    // rom_array[20527] = 32'hFFFFFFF1;
    // rom_array[20528] = 32'hFFFFFFF1;
    // rom_array[20529] = 32'hFFFFFFF0;
    // rom_array[20530] = 32'hFFFFFFF0;
    // rom_array[20531] = 32'hFFFFFFF1;
    // rom_array[20532] = 32'hFFFFFFF1;
    // rom_array[20533] = 32'hFFFFFFF0;
    // rom_array[20534] = 32'hFFFFFFF0;
    // rom_array[20535] = 32'hFFFFFFF1;
    // rom_array[20536] = 32'hFFFFFFF1;
    // rom_array[20537] = 32'hFFFFFFF0;
    // rom_array[20538] = 32'hFFFFFFF0;
    // rom_array[20539] = 32'hFFFFFFF1;
    // rom_array[20540] = 32'hFFFFFFF1;
    // rom_array[20541] = 32'hFFFFFFF0;
    // rom_array[20542] = 32'hFFFFFFF0;
    // rom_array[20543] = 32'hFFFFFFF1;
    // rom_array[20544] = 32'hFFFFFFF1;
    // rom_array[20545] = 32'hFFFFFFF0;
    // rom_array[20546] = 32'hFFFFFFF0;
    // rom_array[20547] = 32'hFFFFFFF1;
    // rom_array[20548] = 32'hFFFFFFF1;
    // rom_array[20549] = 32'hFFFFFFF0;
    // rom_array[20550] = 32'hFFFFFFF0;
    // rom_array[20551] = 32'hFFFFFFF1;
    // rom_array[20552] = 32'hFFFFFFF1;
    // rom_array[20553] = 32'hFFFFFFF0;
    // rom_array[20554] = 32'hFFFFFFF0;
    // rom_array[20555] = 32'hFFFFFFF1;
    // rom_array[20556] = 32'hFFFFFFF1;
    // rom_array[20557] = 32'hFFFFFFF0;
    // rom_array[20558] = 32'hFFFFFFF0;
    // rom_array[20559] = 32'hFFFFFFF1;
    // rom_array[20560] = 32'hFFFFFFF1;
    // rom_array[20561] = 32'hFFFFFFF0;
    // rom_array[20562] = 32'hFFFFFFF0;
    // rom_array[20563] = 32'hFFFFFFF1;
    // rom_array[20564] = 32'hFFFFFFF1;
    // rom_array[20565] = 32'hFFFFFFF0;
    // rom_array[20566] = 32'hFFFFFFF0;
    // rom_array[20567] = 32'hFFFFFFF1;
    // rom_array[20568] = 32'hFFFFFFF1;
    // rom_array[20569] = 32'hFFFFFFF0;
    // rom_array[20570] = 32'hFFFFFFF0;
    // rom_array[20571] = 32'hFFFFFFF1;
    // rom_array[20572] = 32'hFFFFFFF1;
    // rom_array[20573] = 32'hFFFFFFF0;
    // rom_array[20574] = 32'hFFFFFFF0;
    // rom_array[20575] = 32'hFFFFFFF1;
    // rom_array[20576] = 32'hFFFFFFF1;
    // rom_array[20577] = 32'hFFFFFFF0;
    // rom_array[20578] = 32'hFFFFFFF0;
    // rom_array[20579] = 32'hFFFFFFF1;
    // rom_array[20580] = 32'hFFFFFFF1;
    // rom_array[20581] = 32'hFFFFFFF0;
    // rom_array[20582] = 32'hFFFFFFF0;
    // rom_array[20583] = 32'hFFFFFFF1;
    // rom_array[20584] = 32'hFFFFFFF1;
    // rom_array[20585] = 32'hFFFFFFF0;
    // rom_array[20586] = 32'hFFFFFFF0;
    // rom_array[20587] = 32'hFFFFFFF1;
    // rom_array[20588] = 32'hFFFFFFF1;
    // rom_array[20589] = 32'hFFFFFFF0;
    // rom_array[20590] = 32'hFFFFFFF0;
    // rom_array[20591] = 32'hFFFFFFF1;
    // rom_array[20592] = 32'hFFFFFFF1;
    // rom_array[20593] = 32'hFFFFFFF0;
    // rom_array[20594] = 32'hFFFFFFF0;
    // rom_array[20595] = 32'hFFFFFFF1;
    // rom_array[20596] = 32'hFFFFFFF1;
    // rom_array[20597] = 32'hFFFFFFF0;
    // rom_array[20598] = 32'hFFFFFFF0;
    // rom_array[20599] = 32'hFFFFFFF1;
    // rom_array[20600] = 32'hFFFFFFF1;
    // rom_array[20601] = 32'hFFFFFFF1;
    // rom_array[20602] = 32'hFFFFFFF1;
    // rom_array[20603] = 32'hFFFFFFF1;
    // rom_array[20604] = 32'hFFFFFFF1;
    // rom_array[20605] = 32'hFFFFFFF1;
    // rom_array[20606] = 32'hFFFFFFF1;
    // rom_array[20607] = 32'hFFFFFFF1;
    // rom_array[20608] = 32'hFFFFFFF1;
    // rom_array[20609] = 32'hFFFFFFF1;
    // rom_array[20610] = 32'hFFFFFFF1;
    // rom_array[20611] = 32'hFFFFFFF1;
    // rom_array[20612] = 32'hFFFFFFF1;
    // rom_array[20613] = 32'hFFFFFFF1;
    // rom_array[20614] = 32'hFFFFFFF1;
    // rom_array[20615] = 32'hFFFFFFF1;
    // rom_array[20616] = 32'hFFFFFFF1;
    // rom_array[20617] = 32'hFFFFFFF1;
    // rom_array[20618] = 32'hFFFFFFF1;
    // rom_array[20619] = 32'hFFFFFFF1;
    // rom_array[20620] = 32'hFFFFFFF1;
    // rom_array[20621] = 32'hFFFFFFF1;
    // rom_array[20622] = 32'hFFFFFFF1;
    // rom_array[20623] = 32'hFFFFFFF1;
    // rom_array[20624] = 32'hFFFFFFF1;
    // rom_array[20625] = 32'hFFFFFFF1;
    // rom_array[20626] = 32'hFFFFFFF1;
    // rom_array[20627] = 32'hFFFFFFF1;
    // rom_array[20628] = 32'hFFFFFFF1;
    // rom_array[20629] = 32'hFFFFFFF1;
    // rom_array[20630] = 32'hFFFFFFF1;
    // rom_array[20631] = 32'hFFFFFFF1;
    // rom_array[20632] = 32'hFFFFFFF1;
    // rom_array[20633] = 32'hFFFFFFF1;
    // rom_array[20634] = 32'hFFFFFFF1;
    // rom_array[20635] = 32'hFFFFFFF1;
    // rom_array[20636] = 32'hFFFFFFF1;
    // rom_array[20637] = 32'hFFFFFFF1;
    // rom_array[20638] = 32'hFFFFFFF1;
    // rom_array[20639] = 32'hFFFFFFF1;
    // rom_array[20640] = 32'hFFFFFFF1;
    // rom_array[20641] = 32'hFFFFFFF1;
    // rom_array[20642] = 32'hFFFFFFF1;
    // rom_array[20643] = 32'hFFFFFFF1;
    // rom_array[20644] = 32'hFFFFFFF1;
    // rom_array[20645] = 32'hFFFFFFF1;
    // rom_array[20646] = 32'hFFFFFFF1;
    // rom_array[20647] = 32'hFFFFFFF1;
    // rom_array[20648] = 32'hFFFFFFF1;
    // rom_array[20649] = 32'hFFFFFFF1;
    // rom_array[20650] = 32'hFFFFFFF1;
    // rom_array[20651] = 32'hFFFFFFF1;
    // rom_array[20652] = 32'hFFFFFFF1;
    // rom_array[20653] = 32'hFFFFFFF1;
    // rom_array[20654] = 32'hFFFFFFF1;
    // rom_array[20655] = 32'hFFFFFFF1;
    // rom_array[20656] = 32'hFFFFFFF1;
    // rom_array[20657] = 32'hFFFFFFF1;
    // rom_array[20658] = 32'hFFFFFFF1;
    // rom_array[20659] = 32'hFFFFFFF1;
    // rom_array[20660] = 32'hFFFFFFF1;
    // rom_array[20661] = 32'hFFFFFFF1;
    // rom_array[20662] = 32'hFFFFFFF1;
    // rom_array[20663] = 32'hFFFFFFF1;
    // rom_array[20664] = 32'hFFFFFFF1;
    // rom_array[20665] = 32'hFFFFFFF0;
    // rom_array[20666] = 32'hFFFFFFF0;
    // rom_array[20667] = 32'hFFFFFFF1;
    // rom_array[20668] = 32'hFFFFFFF1;
    // rom_array[20669] = 32'hFFFFFFF0;
    // rom_array[20670] = 32'hFFFFFFF0;
    // rom_array[20671] = 32'hFFFFFFF1;
    // rom_array[20672] = 32'hFFFFFFF1;
    // rom_array[20673] = 32'hFFFFFFF0;
    // rom_array[20674] = 32'hFFFFFFF0;
    // rom_array[20675] = 32'hFFFFFFF1;
    // rom_array[20676] = 32'hFFFFFFF1;
    // rom_array[20677] = 32'hFFFFFFF0;
    // rom_array[20678] = 32'hFFFFFFF0;
    // rom_array[20679] = 32'hFFFFFFF1;
    // rom_array[20680] = 32'hFFFFFFF1;
    // rom_array[20681] = 32'hFFFFFFF0;
    // rom_array[20682] = 32'hFFFFFFF0;
    // rom_array[20683] = 32'hFFFFFFF1;
    // rom_array[20684] = 32'hFFFFFFF1;
    // rom_array[20685] = 32'hFFFFFFF0;
    // rom_array[20686] = 32'hFFFFFFF0;
    // rom_array[20687] = 32'hFFFFFFF1;
    // rom_array[20688] = 32'hFFFFFFF1;
    // rom_array[20689] = 32'hFFFFFFF0;
    // rom_array[20690] = 32'hFFFFFFF0;
    // rom_array[20691] = 32'hFFFFFFF1;
    // rom_array[20692] = 32'hFFFFFFF1;
    // rom_array[20693] = 32'hFFFFFFF0;
    // rom_array[20694] = 32'hFFFFFFF0;
    // rom_array[20695] = 32'hFFFFFFF1;
    // rom_array[20696] = 32'hFFFFFFF1;
    // rom_array[20697] = 32'hFFFFFFF0;
    // rom_array[20698] = 32'hFFFFFFF0;
    // rom_array[20699] = 32'hFFFFFFF1;
    // rom_array[20700] = 32'hFFFFFFF1;
    // rom_array[20701] = 32'hFFFFFFF0;
    // rom_array[20702] = 32'hFFFFFFF0;
    // rom_array[20703] = 32'hFFFFFFF1;
    // rom_array[20704] = 32'hFFFFFFF1;
    // rom_array[20705] = 32'hFFFFFFF0;
    // rom_array[20706] = 32'hFFFFFFF0;
    // rom_array[20707] = 32'hFFFFFFF1;
    // rom_array[20708] = 32'hFFFFFFF1;
    // rom_array[20709] = 32'hFFFFFFF0;
    // rom_array[20710] = 32'hFFFFFFF0;
    // rom_array[20711] = 32'hFFFFFFF1;
    // rom_array[20712] = 32'hFFFFFFF1;
    // rom_array[20713] = 32'hFFFFFFF0;
    // rom_array[20714] = 32'hFFFFFFF0;
    // rom_array[20715] = 32'hFFFFFFF1;
    // rom_array[20716] = 32'hFFFFFFF1;
    // rom_array[20717] = 32'hFFFFFFF0;
    // rom_array[20718] = 32'hFFFFFFF0;
    // rom_array[20719] = 32'hFFFFFFF1;
    // rom_array[20720] = 32'hFFFFFFF1;
    // rom_array[20721] = 32'hFFFFFFF0;
    // rom_array[20722] = 32'hFFFFFFF0;
    // rom_array[20723] = 32'hFFFFFFF1;
    // rom_array[20724] = 32'hFFFFFFF1;
    // rom_array[20725] = 32'hFFFFFFF0;
    // rom_array[20726] = 32'hFFFFFFF0;
    // rom_array[20727] = 32'hFFFFFFF1;
    // rom_array[20728] = 32'hFFFFFFF1;
    // rom_array[20729] = 32'hFFFFFFF1;
    // rom_array[20730] = 32'hFFFFFFF1;
    // rom_array[20731] = 32'hFFFFFFF1;
    // rom_array[20732] = 32'hFFFFFFF1;
    // rom_array[20733] = 32'hFFFFFFF1;
    // rom_array[20734] = 32'hFFFFFFF1;
    // rom_array[20735] = 32'hFFFFFFF1;
    // rom_array[20736] = 32'hFFFFFFF1;
    // rom_array[20737] = 32'hFFFFFFF1;
    // rom_array[20738] = 32'hFFFFFFF1;
    // rom_array[20739] = 32'hFFFFFFF1;
    // rom_array[20740] = 32'hFFFFFFF1;
    // rom_array[20741] = 32'hFFFFFFF1;
    // rom_array[20742] = 32'hFFFFFFF1;
    // rom_array[20743] = 32'hFFFFFFF1;
    // rom_array[20744] = 32'hFFFFFFF1;
    // rom_array[20745] = 32'hFFFFFFF1;
    // rom_array[20746] = 32'hFFFFFFF1;
    // rom_array[20747] = 32'hFFFFFFF1;
    // rom_array[20748] = 32'hFFFFFFF1;
    // rom_array[20749] = 32'hFFFFFFF1;
    // rom_array[20750] = 32'hFFFFFFF1;
    // rom_array[20751] = 32'hFFFFFFF1;
    // rom_array[20752] = 32'hFFFFFFF1;
    // rom_array[20753] = 32'hFFFFFFF1;
    // rom_array[20754] = 32'hFFFFFFF1;
    // rom_array[20755] = 32'hFFFFFFF1;
    // rom_array[20756] = 32'hFFFFFFF1;
    // rom_array[20757] = 32'hFFFFFFF1;
    // rom_array[20758] = 32'hFFFFFFF1;
    // rom_array[20759] = 32'hFFFFFFF1;
    // rom_array[20760] = 32'hFFFFFFF1;
    // rom_array[20761] = 32'hFFFFFFF1;
    // rom_array[20762] = 32'hFFFFFFF1;
    // rom_array[20763] = 32'hFFFFFFF1;
    // rom_array[20764] = 32'hFFFFFFF1;
    // rom_array[20765] = 32'hFFFFFFF1;
    // rom_array[20766] = 32'hFFFFFFF1;
    // rom_array[20767] = 32'hFFFFFFF1;
    // rom_array[20768] = 32'hFFFFFFF1;
    // rom_array[20769] = 32'hFFFFFFF1;
    // rom_array[20770] = 32'hFFFFFFF1;
    // rom_array[20771] = 32'hFFFFFFF1;
    // rom_array[20772] = 32'hFFFFFFF1;
    // rom_array[20773] = 32'hFFFFFFF1;
    // rom_array[20774] = 32'hFFFFFFF1;
    // rom_array[20775] = 32'hFFFFFFF1;
    // rom_array[20776] = 32'hFFFFFFF1;
    // rom_array[20777] = 32'hFFFFFFF1;
    // rom_array[20778] = 32'hFFFFFFF1;
    // rom_array[20779] = 32'hFFFFFFF1;
    // rom_array[20780] = 32'hFFFFFFF1;
    // rom_array[20781] = 32'hFFFFFFF1;
    // rom_array[20782] = 32'hFFFFFFF1;
    // rom_array[20783] = 32'hFFFFFFF1;
    // rom_array[20784] = 32'hFFFFFFF1;
    // rom_array[20785] = 32'hFFFFFFF1;
    // rom_array[20786] = 32'hFFFFFFF1;
    // rom_array[20787] = 32'hFFFFFFF1;
    // rom_array[20788] = 32'hFFFFFFF1;
    // rom_array[20789] = 32'hFFFFFFF1;
    // rom_array[20790] = 32'hFFFFFFF1;
    // rom_array[20791] = 32'hFFFFFFF1;
    // rom_array[20792] = 32'hFFFFFFF1;
    // rom_array[20793] = 32'hFFFFFFF0;
    // rom_array[20794] = 32'hFFFFFFF0;
    // rom_array[20795] = 32'hFFFFFFF1;
    // rom_array[20796] = 32'hFFFFFFF1;
    // rom_array[20797] = 32'hFFFFFFF0;
    // rom_array[20798] = 32'hFFFFFFF0;
    // rom_array[20799] = 32'hFFFFFFF1;
    // rom_array[20800] = 32'hFFFFFFF1;
    // rom_array[20801] = 32'hFFFFFFF0;
    // rom_array[20802] = 32'hFFFFFFF0;
    // rom_array[20803] = 32'hFFFFFFF1;
    // rom_array[20804] = 32'hFFFFFFF1;
    // rom_array[20805] = 32'hFFFFFFF0;
    // rom_array[20806] = 32'hFFFFFFF0;
    // rom_array[20807] = 32'hFFFFFFF1;
    // rom_array[20808] = 32'hFFFFFFF1;
    // rom_array[20809] = 32'hFFFFFFF0;
    // rom_array[20810] = 32'hFFFFFFF0;
    // rom_array[20811] = 32'hFFFFFFF1;
    // rom_array[20812] = 32'hFFFFFFF1;
    // rom_array[20813] = 32'hFFFFFFF0;
    // rom_array[20814] = 32'hFFFFFFF0;
    // rom_array[20815] = 32'hFFFFFFF1;
    // rom_array[20816] = 32'hFFFFFFF1;
    // rom_array[20817] = 32'hFFFFFFF0;
    // rom_array[20818] = 32'hFFFFFFF0;
    // rom_array[20819] = 32'hFFFFFFF1;
    // rom_array[20820] = 32'hFFFFFFF1;
    // rom_array[20821] = 32'hFFFFFFF0;
    // rom_array[20822] = 32'hFFFFFFF0;
    // rom_array[20823] = 32'hFFFFFFF1;
    // rom_array[20824] = 32'hFFFFFFF1;
    // rom_array[20825] = 32'hFFFFFFF0;
    // rom_array[20826] = 32'hFFFFFFF0;
    // rom_array[20827] = 32'hFFFFFFF1;
    // rom_array[20828] = 32'hFFFFFFF1;
    // rom_array[20829] = 32'hFFFFFFF0;
    // rom_array[20830] = 32'hFFFFFFF0;
    // rom_array[20831] = 32'hFFFFFFF1;
    // rom_array[20832] = 32'hFFFFFFF1;
    // rom_array[20833] = 32'hFFFFFFF0;
    // rom_array[20834] = 32'hFFFFFFF0;
    // rom_array[20835] = 32'hFFFFFFF1;
    // rom_array[20836] = 32'hFFFFFFF1;
    // rom_array[20837] = 32'hFFFFFFF0;
    // rom_array[20838] = 32'hFFFFFFF0;
    // rom_array[20839] = 32'hFFFFFFF1;
    // rom_array[20840] = 32'hFFFFFFF1;
    // rom_array[20841] = 32'hFFFFFFF0;
    // rom_array[20842] = 32'hFFFFFFF0;
    // rom_array[20843] = 32'hFFFFFFF1;
    // rom_array[20844] = 32'hFFFFFFF1;
    // rom_array[20845] = 32'hFFFFFFF0;
    // rom_array[20846] = 32'hFFFFFFF0;
    // rom_array[20847] = 32'hFFFFFFF1;
    // rom_array[20848] = 32'hFFFFFFF1;
    // rom_array[20849] = 32'hFFFFFFF0;
    // rom_array[20850] = 32'hFFFFFFF0;
    // rom_array[20851] = 32'hFFFFFFF1;
    // rom_array[20852] = 32'hFFFFFFF1;
    // rom_array[20853] = 32'hFFFFFFF0;
    // rom_array[20854] = 32'hFFFFFFF0;
    // rom_array[20855] = 32'hFFFFFFF1;
    // rom_array[20856] = 32'hFFFFFFF1;
    // rom_array[20857] = 32'hFFFFFFF0;
    // rom_array[20858] = 32'hFFFFFFF0;
    // rom_array[20859] = 32'hFFFFFFF0;
    // rom_array[20860] = 32'hFFFFFFF0;
    // rom_array[20861] = 32'hFFFFFFF0;
    // rom_array[20862] = 32'hFFFFFFF0;
    // rom_array[20863] = 32'hFFFFFFF1;
    // rom_array[20864] = 32'hFFFFFFF1;
    // rom_array[20865] = 32'hFFFFFFF0;
    // rom_array[20866] = 32'hFFFFFFF0;
    // rom_array[20867] = 32'hFFFFFFF0;
    // rom_array[20868] = 32'hFFFFFFF0;
    // rom_array[20869] = 32'hFFFFFFF0;
    // rom_array[20870] = 32'hFFFFFFF0;
    // rom_array[20871] = 32'hFFFFFFF1;
    // rom_array[20872] = 32'hFFFFFFF1;
    // rom_array[20873] = 32'hFFFFFFF0;
    // rom_array[20874] = 32'hFFFFFFF0;
    // rom_array[20875] = 32'hFFFFFFF0;
    // rom_array[20876] = 32'hFFFFFFF0;
    // rom_array[20877] = 32'hFFFFFFF1;
    // rom_array[20878] = 32'hFFFFFFF1;
    // rom_array[20879] = 32'hFFFFFFF1;
    // rom_array[20880] = 32'hFFFFFFF1;
    // rom_array[20881] = 32'hFFFFFFF0;
    // rom_array[20882] = 32'hFFFFFFF0;
    // rom_array[20883] = 32'hFFFFFFF0;
    // rom_array[20884] = 32'hFFFFFFF0;
    // rom_array[20885] = 32'hFFFFFFF1;
    // rom_array[20886] = 32'hFFFFFFF1;
    // rom_array[20887] = 32'hFFFFFFF1;
    // rom_array[20888] = 32'hFFFFFFF1;
    // rom_array[20889] = 32'hFFFFFFF0;
    // rom_array[20890] = 32'hFFFFFFF0;
    // rom_array[20891] = 32'hFFFFFFF1;
    // rom_array[20892] = 32'hFFFFFFF1;
    // rom_array[20893] = 32'hFFFFFFF0;
    // rom_array[20894] = 32'hFFFFFFF0;
    // rom_array[20895] = 32'hFFFFFFF1;
    // rom_array[20896] = 32'hFFFFFFF1;
    // rom_array[20897] = 32'hFFFFFFF0;
    // rom_array[20898] = 32'hFFFFFFF0;
    // rom_array[20899] = 32'hFFFFFFF1;
    // rom_array[20900] = 32'hFFFFFFF1;
    // rom_array[20901] = 32'hFFFFFFF0;
    // rom_array[20902] = 32'hFFFFFFF0;
    // rom_array[20903] = 32'hFFFFFFF1;
    // rom_array[20904] = 32'hFFFFFFF1;
    // rom_array[20905] = 32'hFFFFFFF0;
    // rom_array[20906] = 32'hFFFFFFF0;
    // rom_array[20907] = 32'hFFFFFFF1;
    // rom_array[20908] = 32'hFFFFFFF1;
    // rom_array[20909] = 32'hFFFFFFF0;
    // rom_array[20910] = 32'hFFFFFFF0;
    // rom_array[20911] = 32'hFFFFFFF1;
    // rom_array[20912] = 32'hFFFFFFF1;
    // rom_array[20913] = 32'hFFFFFFF0;
    // rom_array[20914] = 32'hFFFFFFF0;
    // rom_array[20915] = 32'hFFFFFFF1;
    // rom_array[20916] = 32'hFFFFFFF1;
    // rom_array[20917] = 32'hFFFFFFF0;
    // rom_array[20918] = 32'hFFFFFFF0;
    // rom_array[20919] = 32'hFFFFFFF1;
    // rom_array[20920] = 32'hFFFFFFF1;
    // rom_array[20921] = 32'hFFFFFFF0;
    // rom_array[20922] = 32'hFFFFFFF0;
    // rom_array[20923] = 32'hFFFFFFF0;
    // rom_array[20924] = 32'hFFFFFFF0;
    // rom_array[20925] = 32'hFFFFFFF1;
    // rom_array[20926] = 32'hFFFFFFF1;
    // rom_array[20927] = 32'hFFFFFFF1;
    // rom_array[20928] = 32'hFFFFFFF1;
    // rom_array[20929] = 32'hFFFFFFF0;
    // rom_array[20930] = 32'hFFFFFFF0;
    // rom_array[20931] = 32'hFFFFFFF0;
    // rom_array[20932] = 32'hFFFFFFF0;
    // rom_array[20933] = 32'hFFFFFFF1;
    // rom_array[20934] = 32'hFFFFFFF1;
    // rom_array[20935] = 32'hFFFFFFF1;
    // rom_array[20936] = 32'hFFFFFFF1;
    // rom_array[20937] = 32'hFFFFFFF0;
    // rom_array[20938] = 32'hFFFFFFF0;
    // rom_array[20939] = 32'hFFFFFFF0;
    // rom_array[20940] = 32'hFFFFFFF0;
    // rom_array[20941] = 32'hFFFFFFF1;
    // rom_array[20942] = 32'hFFFFFFF1;
    // rom_array[20943] = 32'hFFFFFFF1;
    // rom_array[20944] = 32'hFFFFFFF1;
    // rom_array[20945] = 32'hFFFFFFF0;
    // rom_array[20946] = 32'hFFFFFFF0;
    // rom_array[20947] = 32'hFFFFFFF0;
    // rom_array[20948] = 32'hFFFFFFF0;
    // rom_array[20949] = 32'hFFFFFFF1;
    // rom_array[20950] = 32'hFFFFFFF1;
    // rom_array[20951] = 32'hFFFFFFF1;
    // rom_array[20952] = 32'hFFFFFFF1;
    // rom_array[20953] = 32'hFFFFFFF0;
    // rom_array[20954] = 32'hFFFFFFF0;
    // rom_array[20955] = 32'hFFFFFFF0;
    // rom_array[20956] = 32'hFFFFFFF0;
    // rom_array[20957] = 32'hFFFFFFF1;
    // rom_array[20958] = 32'hFFFFFFF1;
    // rom_array[20959] = 32'hFFFFFFF1;
    // rom_array[20960] = 32'hFFFFFFF1;
    // rom_array[20961] = 32'hFFFFFFF0;
    // rom_array[20962] = 32'hFFFFFFF0;
    // rom_array[20963] = 32'hFFFFFFF0;
    // rom_array[20964] = 32'hFFFFFFF0;
    // rom_array[20965] = 32'hFFFFFFF1;
    // rom_array[20966] = 32'hFFFFFFF1;
    // rom_array[20967] = 32'hFFFFFFF1;
    // rom_array[20968] = 32'hFFFFFFF1;
    // rom_array[20969] = 32'hFFFFFFF1;
    // rom_array[20970] = 32'hFFFFFFF1;
    // rom_array[20971] = 32'hFFFFFFF1;
    // rom_array[20972] = 32'hFFFFFFF1;
    // rom_array[20973] = 32'hFFFFFFF1;
    // rom_array[20974] = 32'hFFFFFFF1;
    // rom_array[20975] = 32'hFFFFFFF1;
    // rom_array[20976] = 32'hFFFFFFF1;
    // rom_array[20977] = 32'hFFFFFFF1;
    // rom_array[20978] = 32'hFFFFFFF1;
    // rom_array[20979] = 32'hFFFFFFF1;
    // rom_array[20980] = 32'hFFFFFFF1;
    // rom_array[20981] = 32'hFFFFFFF1;
    // rom_array[20982] = 32'hFFFFFFF1;
    // rom_array[20983] = 32'hFFFFFFF1;
    // rom_array[20984] = 32'hFFFFFFF1;
    // rom_array[20985] = 32'hFFFFFFF1;
    // rom_array[20986] = 32'hFFFFFFF1;
    // rom_array[20987] = 32'hFFFFFFF1;
    // rom_array[20988] = 32'hFFFFFFF1;
    // rom_array[20989] = 32'hFFFFFFF1;
    // rom_array[20990] = 32'hFFFFFFF1;
    // rom_array[20991] = 32'hFFFFFFF1;
    // rom_array[20992] = 32'hFFFFFFF1;
    // rom_array[20993] = 32'hFFFFFFF1;
    // rom_array[20994] = 32'hFFFFFFF1;
    // rom_array[20995] = 32'hFFFFFFF1;
    // rom_array[20996] = 32'hFFFFFFF1;
    // rom_array[20997] = 32'hFFFFFFF1;
    // rom_array[20998] = 32'hFFFFFFF1;
    // rom_array[20999] = 32'hFFFFFFF1;
    // rom_array[21000] = 32'hFFFFFFF1;
    // rom_array[21001] = 32'hFFFFFFF0;
    // rom_array[21002] = 32'hFFFFFFF0;
    // rom_array[21003] = 32'hFFFFFFF0;
    // rom_array[21004] = 32'hFFFFFFF0;
    // rom_array[21005] = 32'hFFFFFFF1;
    // rom_array[21006] = 32'hFFFFFFF1;
    // rom_array[21007] = 32'hFFFFFFF1;
    // rom_array[21008] = 32'hFFFFFFF1;
    // rom_array[21009] = 32'hFFFFFFF0;
    // rom_array[21010] = 32'hFFFFFFF0;
    // rom_array[21011] = 32'hFFFFFFF0;
    // rom_array[21012] = 32'hFFFFFFF0;
    // rom_array[21013] = 32'hFFFFFFF1;
    // rom_array[21014] = 32'hFFFFFFF1;
    // rom_array[21015] = 32'hFFFFFFF1;
    // rom_array[21016] = 32'hFFFFFFF1;
    // rom_array[21017] = 32'hFFFFFFF0;
    // rom_array[21018] = 32'hFFFFFFF0;
    // rom_array[21019] = 32'hFFFFFFF0;
    // rom_array[21020] = 32'hFFFFFFF0;
    // rom_array[21021] = 32'hFFFFFFF1;
    // rom_array[21022] = 32'hFFFFFFF1;
    // rom_array[21023] = 32'hFFFFFFF1;
    // rom_array[21024] = 32'hFFFFFFF1;
    // rom_array[21025] = 32'hFFFFFFF0;
    // rom_array[21026] = 32'hFFFFFFF0;
    // rom_array[21027] = 32'hFFFFFFF0;
    // rom_array[21028] = 32'hFFFFFFF0;
    // rom_array[21029] = 32'hFFFFFFF1;
    // rom_array[21030] = 32'hFFFFFFF1;
    // rom_array[21031] = 32'hFFFFFFF1;
    // rom_array[21032] = 32'hFFFFFFF1;
    // rom_array[21033] = 32'hFFFFFFF0;
    // rom_array[21034] = 32'hFFFFFFF0;
    // rom_array[21035] = 32'hFFFFFFF0;
    // rom_array[21036] = 32'hFFFFFFF0;
    // rom_array[21037] = 32'hFFFFFFF1;
    // rom_array[21038] = 32'hFFFFFFF1;
    // rom_array[21039] = 32'hFFFFFFF1;
    // rom_array[21040] = 32'hFFFFFFF1;
    // rom_array[21041] = 32'hFFFFFFF0;
    // rom_array[21042] = 32'hFFFFFFF0;
    // rom_array[21043] = 32'hFFFFFFF0;
    // rom_array[21044] = 32'hFFFFFFF0;
    // rom_array[21045] = 32'hFFFFFFF1;
    // rom_array[21046] = 32'hFFFFFFF1;
    // rom_array[21047] = 32'hFFFFFFF1;
    // rom_array[21048] = 32'hFFFFFFF1;
    // rom_array[21049] = 32'hFFFFFFF0;
    // rom_array[21050] = 32'hFFFFFFF0;
    // rom_array[21051] = 32'hFFFFFFF0;
    // rom_array[21052] = 32'hFFFFFFF0;
    // rom_array[21053] = 32'hFFFFFFF1;
    // rom_array[21054] = 32'hFFFFFFF1;
    // rom_array[21055] = 32'hFFFFFFF1;
    // rom_array[21056] = 32'hFFFFFFF1;
    // rom_array[21057] = 32'hFFFFFFF0;
    // rom_array[21058] = 32'hFFFFFFF0;
    // rom_array[21059] = 32'hFFFFFFF0;
    // rom_array[21060] = 32'hFFFFFFF0;
    // rom_array[21061] = 32'hFFFFFFF1;
    // rom_array[21062] = 32'hFFFFFFF1;
    // rom_array[21063] = 32'hFFFFFFF1;
    // rom_array[21064] = 32'hFFFFFFF1;
    // rom_array[21065] = 32'hFFFFFFF0;
    // rom_array[21066] = 32'hFFFFFFF0;
    // rom_array[21067] = 32'hFFFFFFF1;
    // rom_array[21068] = 32'hFFFFFFF1;
    // rom_array[21069] = 32'hFFFFFFF0;
    // rom_array[21070] = 32'hFFFFFFF0;
    // rom_array[21071] = 32'hFFFFFFF1;
    // rom_array[21072] = 32'hFFFFFFF1;
    // rom_array[21073] = 32'hFFFFFFF0;
    // rom_array[21074] = 32'hFFFFFFF0;
    // rom_array[21075] = 32'hFFFFFFF1;
    // rom_array[21076] = 32'hFFFFFFF1;
    // rom_array[21077] = 32'hFFFFFFF0;
    // rom_array[21078] = 32'hFFFFFFF0;
    // rom_array[21079] = 32'hFFFFFFF1;
    // rom_array[21080] = 32'hFFFFFFF1;
    // rom_array[21081] = 32'hFFFFFFF0;
    // rom_array[21082] = 32'hFFFFFFF0;
    // rom_array[21083] = 32'hFFFFFFF1;
    // rom_array[21084] = 32'hFFFFFFF1;
    // rom_array[21085] = 32'hFFFFFFF0;
    // rom_array[21086] = 32'hFFFFFFF0;
    // rom_array[21087] = 32'hFFFFFFF1;
    // rom_array[21088] = 32'hFFFFFFF1;
    // rom_array[21089] = 32'hFFFFFFF0;
    // rom_array[21090] = 32'hFFFFFFF0;
    // rom_array[21091] = 32'hFFFFFFF1;
    // rom_array[21092] = 32'hFFFFFFF1;
    // rom_array[21093] = 32'hFFFFFFF0;
    // rom_array[21094] = 32'hFFFFFFF0;
    // rom_array[21095] = 32'hFFFFFFF1;
    // rom_array[21096] = 32'hFFFFFFF1;
    // rom_array[21097] = 32'hFFFFFFF0;
    // rom_array[21098] = 32'hFFFFFFF0;
    // rom_array[21099] = 32'hFFFFFFF0;
    // rom_array[21100] = 32'hFFFFFFF0;
    // rom_array[21101] = 32'hFFFFFFF1;
    // rom_array[21102] = 32'hFFFFFFF1;
    // rom_array[21103] = 32'hFFFFFFF1;
    // rom_array[21104] = 32'hFFFFFFF1;
    // rom_array[21105] = 32'hFFFFFFF0;
    // rom_array[21106] = 32'hFFFFFFF0;
    // rom_array[21107] = 32'hFFFFFFF0;
    // rom_array[21108] = 32'hFFFFFFF0;
    // rom_array[21109] = 32'hFFFFFFF1;
    // rom_array[21110] = 32'hFFFFFFF1;
    // rom_array[21111] = 32'hFFFFFFF1;
    // rom_array[21112] = 32'hFFFFFFF1;
    // rom_array[21113] = 32'hFFFFFFF0;
    // rom_array[21114] = 32'hFFFFFFF0;
    // rom_array[21115] = 32'hFFFFFFF0;
    // rom_array[21116] = 32'hFFFFFFF0;
    // rom_array[21117] = 32'hFFFFFFF1;
    // rom_array[21118] = 32'hFFFFFFF1;
    // rom_array[21119] = 32'hFFFFFFF1;
    // rom_array[21120] = 32'hFFFFFFF1;
    // rom_array[21121] = 32'hFFFFFFF0;
    // rom_array[21122] = 32'hFFFFFFF0;
    // rom_array[21123] = 32'hFFFFFFF0;
    // rom_array[21124] = 32'hFFFFFFF0;
    // rom_array[21125] = 32'hFFFFFFF1;
    // rom_array[21126] = 32'hFFFFFFF1;
    // rom_array[21127] = 32'hFFFFFFF1;
    // rom_array[21128] = 32'hFFFFFFF1;
    // rom_array[21129] = 32'hFFFFFFF0;
    // rom_array[21130] = 32'hFFFFFFF0;
    // rom_array[21131] = 32'hFFFFFFF1;
    // rom_array[21132] = 32'hFFFFFFF1;
    // rom_array[21133] = 32'hFFFFFFF1;
    // rom_array[21134] = 32'hFFFFFFF1;
    // rom_array[21135] = 32'hFFFFFFF1;
    // rom_array[21136] = 32'hFFFFFFF1;
    // rom_array[21137] = 32'hFFFFFFF0;
    // rom_array[21138] = 32'hFFFFFFF0;
    // rom_array[21139] = 32'hFFFFFFF1;
    // rom_array[21140] = 32'hFFFFFFF1;
    // rom_array[21141] = 32'hFFFFFFF1;
    // rom_array[21142] = 32'hFFFFFFF1;
    // rom_array[21143] = 32'hFFFFFFF1;
    // rom_array[21144] = 32'hFFFFFFF1;
    // rom_array[21145] = 32'hFFFFFFF1;
    // rom_array[21146] = 32'hFFFFFFF1;
    // rom_array[21147] = 32'hFFFFFFF1;
    // rom_array[21148] = 32'hFFFFFFF1;
    // rom_array[21149] = 32'hFFFFFFF1;
    // rom_array[21150] = 32'hFFFFFFF1;
    // rom_array[21151] = 32'hFFFFFFF1;
    // rom_array[21152] = 32'hFFFFFFF1;
    // rom_array[21153] = 32'hFFFFFFF1;
    // rom_array[21154] = 32'hFFFFFFF1;
    // rom_array[21155] = 32'hFFFFFFF1;
    // rom_array[21156] = 32'hFFFFFFF1;
    // rom_array[21157] = 32'hFFFFFFF1;
    // rom_array[21158] = 32'hFFFFFFF1;
    // rom_array[21159] = 32'hFFFFFFF1;
    // rom_array[21160] = 32'hFFFFFFF1;
    // rom_array[21161] = 32'hFFFFFFF1;
    // rom_array[21162] = 32'hFFFFFFF1;
    // rom_array[21163] = 32'hFFFFFFF1;
    // rom_array[21164] = 32'hFFFFFFF1;
    // rom_array[21165] = 32'hFFFFFFF0;
    // rom_array[21166] = 32'hFFFFFFF0;
    // rom_array[21167] = 32'hFFFFFFF0;
    // rom_array[21168] = 32'hFFFFFFF0;
    // rom_array[21169] = 32'hFFFFFFF1;
    // rom_array[21170] = 32'hFFFFFFF1;
    // rom_array[21171] = 32'hFFFFFFF1;
    // rom_array[21172] = 32'hFFFFFFF1;
    // rom_array[21173] = 32'hFFFFFFF0;
    // rom_array[21174] = 32'hFFFFFFF0;
    // rom_array[21175] = 32'hFFFFFFF0;
    // rom_array[21176] = 32'hFFFFFFF0;
    // rom_array[21177] = 32'hFFFFFFF1;
    // rom_array[21178] = 32'hFFFFFFF1;
    // rom_array[21179] = 32'hFFFFFFF1;
    // rom_array[21180] = 32'hFFFFFFF1;
    // rom_array[21181] = 32'hFFFFFFF0;
    // rom_array[21182] = 32'hFFFFFFF0;
    // rom_array[21183] = 32'hFFFFFFF0;
    // rom_array[21184] = 32'hFFFFFFF0;
    // rom_array[21185] = 32'hFFFFFFF1;
    // rom_array[21186] = 32'hFFFFFFF1;
    // rom_array[21187] = 32'hFFFFFFF1;
    // rom_array[21188] = 32'hFFFFFFF1;
    // rom_array[21189] = 32'hFFFFFFF0;
    // rom_array[21190] = 32'hFFFFFFF0;
    // rom_array[21191] = 32'hFFFFFFF0;
    // rom_array[21192] = 32'hFFFFFFF0;
    // rom_array[21193] = 32'hFFFFFFF1;
    // rom_array[21194] = 32'hFFFFFFF1;
    // rom_array[21195] = 32'hFFFFFFF1;
    // rom_array[21196] = 32'hFFFFFFF1;
    // rom_array[21197] = 32'hFFFFFFF0;
    // rom_array[21198] = 32'hFFFFFFF0;
    // rom_array[21199] = 32'hFFFFFFF0;
    // rom_array[21200] = 32'hFFFFFFF0;
    // rom_array[21201] = 32'hFFFFFFF1;
    // rom_array[21202] = 32'hFFFFFFF1;
    // rom_array[21203] = 32'hFFFFFFF1;
    // rom_array[21204] = 32'hFFFFFFF1;
    // rom_array[21205] = 32'hFFFFFFF0;
    // rom_array[21206] = 32'hFFFFFFF0;
    // rom_array[21207] = 32'hFFFFFFF0;
    // rom_array[21208] = 32'hFFFFFFF0;
    // rom_array[21209] = 32'hFFFFFFF1;
    // rom_array[21210] = 32'hFFFFFFF1;
    // rom_array[21211] = 32'hFFFFFFF1;
    // rom_array[21212] = 32'hFFFFFFF1;
    // rom_array[21213] = 32'hFFFFFFF0;
    // rom_array[21214] = 32'hFFFFFFF0;
    // rom_array[21215] = 32'hFFFFFFF0;
    // rom_array[21216] = 32'hFFFFFFF0;
    // rom_array[21217] = 32'hFFFFFFF1;
    // rom_array[21218] = 32'hFFFFFFF1;
    // rom_array[21219] = 32'hFFFFFFF1;
    // rom_array[21220] = 32'hFFFFFFF1;
    // rom_array[21221] = 32'hFFFFFFF0;
    // rom_array[21222] = 32'hFFFFFFF0;
    // rom_array[21223] = 32'hFFFFFFF0;
    // rom_array[21224] = 32'hFFFFFFF0;
    // rom_array[21225] = 32'hFFFFFFF1;
    // rom_array[21226] = 32'hFFFFFFF1;
    // rom_array[21227] = 32'hFFFFFFF1;
    // rom_array[21228] = 32'hFFFFFFF1;
    // rom_array[21229] = 32'hFFFFFFF1;
    // rom_array[21230] = 32'hFFFFFFF1;
    // rom_array[21231] = 32'hFFFFFFF1;
    // rom_array[21232] = 32'hFFFFFFF1;
    // rom_array[21233] = 32'hFFFFFFF1;
    // rom_array[21234] = 32'hFFFFFFF1;
    // rom_array[21235] = 32'hFFFFFFF1;
    // rom_array[21236] = 32'hFFFFFFF1;
    // rom_array[21237] = 32'hFFFFFFF1;
    // rom_array[21238] = 32'hFFFFFFF1;
    // rom_array[21239] = 32'hFFFFFFF1;
    // rom_array[21240] = 32'hFFFFFFF1;
    // rom_array[21241] = 32'hFFFFFFF1;
    // rom_array[21242] = 32'hFFFFFFF1;
    // rom_array[21243] = 32'hFFFFFFF1;
    // rom_array[21244] = 32'hFFFFFFF1;
    // rom_array[21245] = 32'hFFFFFFF1;
    // rom_array[21246] = 32'hFFFFFFF1;
    // rom_array[21247] = 32'hFFFFFFF1;
    // rom_array[21248] = 32'hFFFFFFF1;
    // rom_array[21249] = 32'hFFFFFFF1;
    // rom_array[21250] = 32'hFFFFFFF1;
    // rom_array[21251] = 32'hFFFFFFF1;
    // rom_array[21252] = 32'hFFFFFFF1;
    // rom_array[21253] = 32'hFFFFFFF1;
    // rom_array[21254] = 32'hFFFFFFF1;
    // rom_array[21255] = 32'hFFFFFFF1;
    // rom_array[21256] = 32'hFFFFFFF1;
    // rom_array[21257] = 32'hFFFFFFF1;
    // rom_array[21258] = 32'hFFFFFFF1;
    // rom_array[21259] = 32'hFFFFFFF1;
    // rom_array[21260] = 32'hFFFFFFF1;
    // rom_array[21261] = 32'hFFFFFFF0;
    // rom_array[21262] = 32'hFFFFFFF0;
    // rom_array[21263] = 32'hFFFFFFF0;
    // rom_array[21264] = 32'hFFFFFFF0;
    // rom_array[21265] = 32'hFFFFFFF1;
    // rom_array[21266] = 32'hFFFFFFF1;
    // rom_array[21267] = 32'hFFFFFFF1;
    // rom_array[21268] = 32'hFFFFFFF1;
    // rom_array[21269] = 32'hFFFFFFF0;
    // rom_array[21270] = 32'hFFFFFFF0;
    // rom_array[21271] = 32'hFFFFFFF0;
    // rom_array[21272] = 32'hFFFFFFF0;
    // rom_array[21273] = 32'hFFFFFFF1;
    // rom_array[21274] = 32'hFFFFFFF1;
    // rom_array[21275] = 32'hFFFFFFF1;
    // rom_array[21276] = 32'hFFFFFFF1;
    // rom_array[21277] = 32'hFFFFFFF0;
    // rom_array[21278] = 32'hFFFFFFF0;
    // rom_array[21279] = 32'hFFFFFFF0;
    // rom_array[21280] = 32'hFFFFFFF0;
    // rom_array[21281] = 32'hFFFFFFF1;
    // rom_array[21282] = 32'hFFFFFFF1;
    // rom_array[21283] = 32'hFFFFFFF1;
    // rom_array[21284] = 32'hFFFFFFF1;
    // rom_array[21285] = 32'hFFFFFFF0;
    // rom_array[21286] = 32'hFFFFFFF0;
    // rom_array[21287] = 32'hFFFFFFF0;
    // rom_array[21288] = 32'hFFFFFFF0;
    // rom_array[21289] = 32'hFFFFFFF1;
    // rom_array[21290] = 32'hFFFFFFF1;
    // rom_array[21291] = 32'hFFFFFFF1;
    // rom_array[21292] = 32'hFFFFFFF1;
    // rom_array[21293] = 32'hFFFFFFF0;
    // rom_array[21294] = 32'hFFFFFFF0;
    // rom_array[21295] = 32'hFFFFFFF1;
    // rom_array[21296] = 32'hFFFFFFF1;
    // rom_array[21297] = 32'hFFFFFFF1;
    // rom_array[21298] = 32'hFFFFFFF1;
    // rom_array[21299] = 32'hFFFFFFF1;
    // rom_array[21300] = 32'hFFFFFFF1;
    // rom_array[21301] = 32'hFFFFFFF0;
    // rom_array[21302] = 32'hFFFFFFF0;
    // rom_array[21303] = 32'hFFFFFFF1;
    // rom_array[21304] = 32'hFFFFFFF1;
    // rom_array[21305] = 32'hFFFFFFF0;
    // rom_array[21306] = 32'hFFFFFFF0;
    // rom_array[21307] = 32'hFFFFFFF1;
    // rom_array[21308] = 32'hFFFFFFF1;
    // rom_array[21309] = 32'hFFFFFFF0;
    // rom_array[21310] = 32'hFFFFFFF0;
    // rom_array[21311] = 32'hFFFFFFF1;
    // rom_array[21312] = 32'hFFFFFFF1;
    // rom_array[21313] = 32'hFFFFFFF0;
    // rom_array[21314] = 32'hFFFFFFF0;
    // rom_array[21315] = 32'hFFFFFFF1;
    // rom_array[21316] = 32'hFFFFFFF1;
    // rom_array[21317] = 32'hFFFFFFF0;
    // rom_array[21318] = 32'hFFFFFFF0;
    // rom_array[21319] = 32'hFFFFFFF1;
    // rom_array[21320] = 32'hFFFFFFF1;
    // rom_array[21321] = 32'hFFFFFFF1;
    // rom_array[21322] = 32'hFFFFFFF1;
    // rom_array[21323] = 32'hFFFFFFF1;
    // rom_array[21324] = 32'hFFFFFFF1;
    // rom_array[21325] = 32'hFFFFFFF1;
    // rom_array[21326] = 32'hFFFFFFF1;
    // rom_array[21327] = 32'hFFFFFFF1;
    // rom_array[21328] = 32'hFFFFFFF1;
    // rom_array[21329] = 32'hFFFFFFF1;
    // rom_array[21330] = 32'hFFFFFFF1;
    // rom_array[21331] = 32'hFFFFFFF1;
    // rom_array[21332] = 32'hFFFFFFF1;
    // rom_array[21333] = 32'hFFFFFFF1;
    // rom_array[21334] = 32'hFFFFFFF1;
    // rom_array[21335] = 32'hFFFFFFF1;
    // rom_array[21336] = 32'hFFFFFFF1;
    // rom_array[21337] = 32'hFFFFFFF1;
    // rom_array[21338] = 32'hFFFFFFF1;
    // rom_array[21339] = 32'hFFFFFFF1;
    // rom_array[21340] = 32'hFFFFFFF1;
    // rom_array[21341] = 32'hFFFFFFF1;
    // rom_array[21342] = 32'hFFFFFFF1;
    // rom_array[21343] = 32'hFFFFFFF1;
    // rom_array[21344] = 32'hFFFFFFF1;
    // rom_array[21345] = 32'hFFFFFFF1;
    // rom_array[21346] = 32'hFFFFFFF1;
    // rom_array[21347] = 32'hFFFFFFF1;
    // rom_array[21348] = 32'hFFFFFFF1;
    // rom_array[21349] = 32'hFFFFFFF1;
    // rom_array[21350] = 32'hFFFFFFF1;
    // rom_array[21351] = 32'hFFFFFFF1;
    // rom_array[21352] = 32'hFFFFFFF1;
    // rom_array[21353] = 32'hFFFFFFF1;
    // rom_array[21354] = 32'hFFFFFFF1;
    // rom_array[21355] = 32'hFFFFFFF1;
    // rom_array[21356] = 32'hFFFFFFF1;
    // rom_array[21357] = 32'hFFFFFFF1;
    // rom_array[21358] = 32'hFFFFFFF1;
    // rom_array[21359] = 32'hFFFFFFF1;
    // rom_array[21360] = 32'hFFFFFFF1;
    // rom_array[21361] = 32'hFFFFFFF1;
    // rom_array[21362] = 32'hFFFFFFF1;
    // rom_array[21363] = 32'hFFFFFFF1;
    // rom_array[21364] = 32'hFFFFFFF1;
    // rom_array[21365] = 32'hFFFFFFF1;
    // rom_array[21366] = 32'hFFFFFFF1;
    // rom_array[21367] = 32'hFFFFFFF1;
    // rom_array[21368] = 32'hFFFFFFF1;
    // rom_array[21369] = 32'hFFFFFFF1;
    // rom_array[21370] = 32'hFFFFFFF1;
    // rom_array[21371] = 32'hFFFFFFF1;
    // rom_array[21372] = 32'hFFFFFFF1;
    // rom_array[21373] = 32'hFFFFFFF1;
    // rom_array[21374] = 32'hFFFFFFF1;
    // rom_array[21375] = 32'hFFFFFFF1;
    // rom_array[21376] = 32'hFFFFFFF1;
    // rom_array[21377] = 32'hFFFFFFF1;
    // rom_array[21378] = 32'hFFFFFFF1;
    // rom_array[21379] = 32'hFFFFFFF1;
    // rom_array[21380] = 32'hFFFFFFF1;
    // rom_array[21381] = 32'hFFFFFFF1;
    // rom_array[21382] = 32'hFFFFFFF1;
    // rom_array[21383] = 32'hFFFFFFF1;
    // rom_array[21384] = 32'hFFFFFFF1;
    // rom_array[21385] = 32'hFFFFFFF1;
    // rom_array[21386] = 32'hFFFFFFF1;
    // rom_array[21387] = 32'hFFFFFFF1;
    // rom_array[21388] = 32'hFFFFFFF1;
    // rom_array[21389] = 32'hFFFFFFF1;
    // rom_array[21390] = 32'hFFFFFFF1;
    // rom_array[21391] = 32'hFFFFFFF1;
    // rom_array[21392] = 32'hFFFFFFF1;
    // rom_array[21393] = 32'hFFFFFFF1;
    // rom_array[21394] = 32'hFFFFFFF1;
    // rom_array[21395] = 32'hFFFFFFF1;
    // rom_array[21396] = 32'hFFFFFFF1;
    // rom_array[21397] = 32'hFFFFFFF1;
    // rom_array[21398] = 32'hFFFFFFF1;
    // rom_array[21399] = 32'hFFFFFFF1;
    // rom_array[21400] = 32'hFFFFFFF1;
    // rom_array[21401] = 32'hFFFFFFF1;
    // rom_array[21402] = 32'hFFFFFFF1;
    // rom_array[21403] = 32'hFFFFFFF1;
    // rom_array[21404] = 32'hFFFFFFF1;
    // rom_array[21405] = 32'hFFFFFFF1;
    // rom_array[21406] = 32'hFFFFFFF1;
    // rom_array[21407] = 32'hFFFFFFF1;
    // rom_array[21408] = 32'hFFFFFFF1;
    // rom_array[21409] = 32'hFFFFFFF1;
    // rom_array[21410] = 32'hFFFFFFF1;
    // rom_array[21411] = 32'hFFFFFFF1;
    // rom_array[21412] = 32'hFFFFFFF1;
    // rom_array[21413] = 32'hFFFFFFF1;
    // rom_array[21414] = 32'hFFFFFFF1;
    // rom_array[21415] = 32'hFFFFFFF1;
    // rom_array[21416] = 32'hFFFFFFF1;
    // rom_array[21417] = 32'hFFFFFFF1;
    // rom_array[21418] = 32'hFFFFFFF1;
    // rom_array[21419] = 32'hFFFFFFF1;
    // rom_array[21420] = 32'hFFFFFFF1;
    // rom_array[21421] = 32'hFFFFFFF1;
    // rom_array[21422] = 32'hFFFFFFF1;
    // rom_array[21423] = 32'hFFFFFFF1;
    // rom_array[21424] = 32'hFFFFFFF1;
    // rom_array[21425] = 32'hFFFFFFF1;
    // rom_array[21426] = 32'hFFFFFFF1;
    // rom_array[21427] = 32'hFFFFFFF1;
    // rom_array[21428] = 32'hFFFFFFF1;
    // rom_array[21429] = 32'hFFFFFFF1;
    // rom_array[21430] = 32'hFFFFFFF1;
    // rom_array[21431] = 32'hFFFFFFF1;
    // rom_array[21432] = 32'hFFFFFFF1;
    // rom_array[21433] = 32'hFFFFFFF1;
    // rom_array[21434] = 32'hFFFFFFF1;
    // rom_array[21435] = 32'hFFFFFFF1;
    // rom_array[21436] = 32'hFFFFFFF1;
    // rom_array[21437] = 32'hFFFFFFF1;
    // rom_array[21438] = 32'hFFFFFFF1;
    // rom_array[21439] = 32'hFFFFFFF1;
    // rom_array[21440] = 32'hFFFFFFF1;
    // rom_array[21441] = 32'hFFFFFFF1;
    // rom_array[21442] = 32'hFFFFFFF1;
    // rom_array[21443] = 32'hFFFFFFF1;
    // rom_array[21444] = 32'hFFFFFFF1;
    // rom_array[21445] = 32'hFFFFFFF1;
    // rom_array[21446] = 32'hFFFFFFF1;
    // rom_array[21447] = 32'hFFFFFFF1;
    // rom_array[21448] = 32'hFFFFFFF1;
    // rom_array[21449] = 32'hFFFFFFF0;
    // rom_array[21450] = 32'hFFFFFFF0;
    // rom_array[21451] = 32'hFFFFFFF1;
    // rom_array[21452] = 32'hFFFFFFF1;
    // rom_array[21453] = 32'hFFFFFFF0;
    // rom_array[21454] = 32'hFFFFFFF0;
    // rom_array[21455] = 32'hFFFFFFF1;
    // rom_array[21456] = 32'hFFFFFFF1;
    // rom_array[21457] = 32'hFFFFFFF0;
    // rom_array[21458] = 32'hFFFFFFF0;
    // rom_array[21459] = 32'hFFFFFFF1;
    // rom_array[21460] = 32'hFFFFFFF1;
    // rom_array[21461] = 32'hFFFFFFF0;
    // rom_array[21462] = 32'hFFFFFFF0;
    // rom_array[21463] = 32'hFFFFFFF1;
    // rom_array[21464] = 32'hFFFFFFF1;
    // rom_array[21465] = 32'hFFFFFFF0;
    // rom_array[21466] = 32'hFFFFFFF0;
    // rom_array[21467] = 32'hFFFFFFF1;
    // rom_array[21468] = 32'hFFFFFFF1;
    // rom_array[21469] = 32'hFFFFFFF0;
    // rom_array[21470] = 32'hFFFFFFF0;
    // rom_array[21471] = 32'hFFFFFFF1;
    // rom_array[21472] = 32'hFFFFFFF1;
    // rom_array[21473] = 32'hFFFFFFF0;
    // rom_array[21474] = 32'hFFFFFFF0;
    // rom_array[21475] = 32'hFFFFFFF1;
    // rom_array[21476] = 32'hFFFFFFF1;
    // rom_array[21477] = 32'hFFFFFFF0;
    // rom_array[21478] = 32'hFFFFFFF0;
    // rom_array[21479] = 32'hFFFFFFF1;
    // rom_array[21480] = 32'hFFFFFFF1;
    // rom_array[21481] = 32'hFFFFFFF0;
    // rom_array[21482] = 32'hFFFFFFF0;
    // rom_array[21483] = 32'hFFFFFFF1;
    // rom_array[21484] = 32'hFFFFFFF1;
    // rom_array[21485] = 32'hFFFFFFF0;
    // rom_array[21486] = 32'hFFFFFFF0;
    // rom_array[21487] = 32'hFFFFFFF1;
    // rom_array[21488] = 32'hFFFFFFF1;
    // rom_array[21489] = 32'hFFFFFFF0;
    // rom_array[21490] = 32'hFFFFFFF0;
    // rom_array[21491] = 32'hFFFFFFF1;
    // rom_array[21492] = 32'hFFFFFFF1;
    // rom_array[21493] = 32'hFFFFFFF0;
    // rom_array[21494] = 32'hFFFFFFF0;
    // rom_array[21495] = 32'hFFFFFFF1;
    // rom_array[21496] = 32'hFFFFFFF1;
    // rom_array[21497] = 32'hFFFFFFF0;
    // rom_array[21498] = 32'hFFFFFFF0;
    // rom_array[21499] = 32'hFFFFFFF1;
    // rom_array[21500] = 32'hFFFFFFF1;
    // rom_array[21501] = 32'hFFFFFFF0;
    // rom_array[21502] = 32'hFFFFFFF0;
    // rom_array[21503] = 32'hFFFFFFF0;
    // rom_array[21504] = 32'hFFFFFFF0;
    // rom_array[21505] = 32'hFFFFFFF0;
    // rom_array[21506] = 32'hFFFFFFF0;
    // rom_array[21507] = 32'hFFFFFFF1;
    // rom_array[21508] = 32'hFFFFFFF1;
    // rom_array[21509] = 32'hFFFFFFF0;
    // rom_array[21510] = 32'hFFFFFFF0;
    // rom_array[21511] = 32'hFFFFFFF0;
    // rom_array[21512] = 32'hFFFFFFF0;
    // rom_array[21513] = 32'hFFFFFFF1;
    // rom_array[21514] = 32'hFFFFFFF1;
    // rom_array[21515] = 32'hFFFFFFF1;
    // rom_array[21516] = 32'hFFFFFFF1;
    // rom_array[21517] = 32'hFFFFFFF0;
    // rom_array[21518] = 32'hFFFFFFF0;
    // rom_array[21519] = 32'hFFFFFFF0;
    // rom_array[21520] = 32'hFFFFFFF0;
    // rom_array[21521] = 32'hFFFFFFF1;
    // rom_array[21522] = 32'hFFFFFFF1;
    // rom_array[21523] = 32'hFFFFFFF1;
    // rom_array[21524] = 32'hFFFFFFF1;
    // rom_array[21525] = 32'hFFFFFFF0;
    // rom_array[21526] = 32'hFFFFFFF0;
    // rom_array[21527] = 32'hFFFFFFF0;
    // rom_array[21528] = 32'hFFFFFFF0;
    // rom_array[21529] = 32'hFFFFFFF1;
    // rom_array[21530] = 32'hFFFFFFF1;
    // rom_array[21531] = 32'hFFFFFFF1;
    // rom_array[21532] = 32'hFFFFFFF1;
    // rom_array[21533] = 32'hFFFFFFF1;
    // rom_array[21534] = 32'hFFFFFFF1;
    // rom_array[21535] = 32'hFFFFFFF1;
    // rom_array[21536] = 32'hFFFFFFF1;
    // rom_array[21537] = 32'hFFFFFFF1;
    // rom_array[21538] = 32'hFFFFFFF1;
    // rom_array[21539] = 32'hFFFFFFF1;
    // rom_array[21540] = 32'hFFFFFFF1;
    // rom_array[21541] = 32'hFFFFFFF1;
    // rom_array[21542] = 32'hFFFFFFF1;
    // rom_array[21543] = 32'hFFFFFFF1;
    // rom_array[21544] = 32'hFFFFFFF1;
    // rom_array[21545] = 32'hFFFFFFF1;
    // rom_array[21546] = 32'hFFFFFFF1;
    // rom_array[21547] = 32'hFFFFFFF1;
    // rom_array[21548] = 32'hFFFFFFF1;
    // rom_array[21549] = 32'hFFFFFFF1;
    // rom_array[21550] = 32'hFFFFFFF1;
    // rom_array[21551] = 32'hFFFFFFF1;
    // rom_array[21552] = 32'hFFFFFFF1;
    // rom_array[21553] = 32'hFFFFFFF1;
    // rom_array[21554] = 32'hFFFFFFF1;
    // rom_array[21555] = 32'hFFFFFFF1;
    // rom_array[21556] = 32'hFFFFFFF1;
    // rom_array[21557] = 32'hFFFFFFF1;
    // rom_array[21558] = 32'hFFFFFFF1;
    // rom_array[21559] = 32'hFFFFFFF1;
    // rom_array[21560] = 32'hFFFFFFF1;
    // rom_array[21561] = 32'hFFFFFFF1;
    // rom_array[21562] = 32'hFFFFFFF1;
    // rom_array[21563] = 32'hFFFFFFF1;
    // rom_array[21564] = 32'hFFFFFFF1;
    // rom_array[21565] = 32'hFFFFFFF0;
    // rom_array[21566] = 32'hFFFFFFF0;
    // rom_array[21567] = 32'hFFFFFFF0;
    // rom_array[21568] = 32'hFFFFFFF0;
    // rom_array[21569] = 32'hFFFFFFF1;
    // rom_array[21570] = 32'hFFFFFFF1;
    // rom_array[21571] = 32'hFFFFFFF1;
    // rom_array[21572] = 32'hFFFFFFF1;
    // rom_array[21573] = 32'hFFFFFFF0;
    // rom_array[21574] = 32'hFFFFFFF0;
    // rom_array[21575] = 32'hFFFFFFF0;
    // rom_array[21576] = 32'hFFFFFFF0;
    // rom_array[21577] = 32'hFFFFFFF1;
    // rom_array[21578] = 32'hFFFFFFF1;
    // rom_array[21579] = 32'hFFFFFFF1;
    // rom_array[21580] = 32'hFFFFFFF1;
    // rom_array[21581] = 32'hFFFFFFF0;
    // rom_array[21582] = 32'hFFFFFFF0;
    // rom_array[21583] = 32'hFFFFFFF0;
    // rom_array[21584] = 32'hFFFFFFF0;
    // rom_array[21585] = 32'hFFFFFFF1;
    // rom_array[21586] = 32'hFFFFFFF1;
    // rom_array[21587] = 32'hFFFFFFF1;
    // rom_array[21588] = 32'hFFFFFFF1;
    // rom_array[21589] = 32'hFFFFFFF0;
    // rom_array[21590] = 32'hFFFFFFF0;
    // rom_array[21591] = 32'hFFFFFFF0;
    // rom_array[21592] = 32'hFFFFFFF0;
    // rom_array[21593] = 32'hFFFFFFF1;
    // rom_array[21594] = 32'hFFFFFFF1;
    // rom_array[21595] = 32'hFFFFFFF1;
    // rom_array[21596] = 32'hFFFFFFF1;
    // rom_array[21597] = 32'hFFFFFFF1;
    // rom_array[21598] = 32'hFFFFFFF1;
    // rom_array[21599] = 32'hFFFFFFF1;
    // rom_array[21600] = 32'hFFFFFFF1;
    // rom_array[21601] = 32'hFFFFFFF1;
    // rom_array[21602] = 32'hFFFFFFF1;
    // rom_array[21603] = 32'hFFFFFFF1;
    // rom_array[21604] = 32'hFFFFFFF1;
    // rom_array[21605] = 32'hFFFFFFF1;
    // rom_array[21606] = 32'hFFFFFFF1;
    // rom_array[21607] = 32'hFFFFFFF1;
    // rom_array[21608] = 32'hFFFFFFF1;
    // rom_array[21609] = 32'hFFFFFFF1;
    // rom_array[21610] = 32'hFFFFFFF1;
    // rom_array[21611] = 32'hFFFFFFF1;
    // rom_array[21612] = 32'hFFFFFFF1;
    // rom_array[21613] = 32'hFFFFFFF0;
    // rom_array[21614] = 32'hFFFFFFF0;
    // rom_array[21615] = 32'hFFFFFFF0;
    // rom_array[21616] = 32'hFFFFFFF0;
    // rom_array[21617] = 32'hFFFFFFF1;
    // rom_array[21618] = 32'hFFFFFFF1;
    // rom_array[21619] = 32'hFFFFFFF1;
    // rom_array[21620] = 32'hFFFFFFF1;
    // rom_array[21621] = 32'hFFFFFFF0;
    // rom_array[21622] = 32'hFFFFFFF0;
    // rom_array[21623] = 32'hFFFFFFF0;
    // rom_array[21624] = 32'hFFFFFFF0;
    // rom_array[21625] = 32'hFFFFFFF0;
    // rom_array[21626] = 32'hFFFFFFF0;
    // rom_array[21627] = 32'hFFFFFFF0;
    // rom_array[21628] = 32'hFFFFFFF0;
    // rom_array[21629] = 32'hFFFFFFF1;
    // rom_array[21630] = 32'hFFFFFFF1;
    // rom_array[21631] = 32'hFFFFFFF1;
    // rom_array[21632] = 32'hFFFFFFF1;
    // rom_array[21633] = 32'hFFFFFFF0;
    // rom_array[21634] = 32'hFFFFFFF0;
    // rom_array[21635] = 32'hFFFFFFF0;
    // rom_array[21636] = 32'hFFFFFFF0;
    // rom_array[21637] = 32'hFFFFFFF1;
    // rom_array[21638] = 32'hFFFFFFF1;
    // rom_array[21639] = 32'hFFFFFFF1;
    // rom_array[21640] = 32'hFFFFFFF1;
    // rom_array[21641] = 32'hFFFFFFF0;
    // rom_array[21642] = 32'hFFFFFFF0;
    // rom_array[21643] = 32'hFFFFFFF0;
    // rom_array[21644] = 32'hFFFFFFF0;
    // rom_array[21645] = 32'hFFFFFFF1;
    // rom_array[21646] = 32'hFFFFFFF1;
    // rom_array[21647] = 32'hFFFFFFF1;
    // rom_array[21648] = 32'hFFFFFFF1;
    // rom_array[21649] = 32'hFFFFFFF0;
    // rom_array[21650] = 32'hFFFFFFF0;
    // rom_array[21651] = 32'hFFFFFFF0;
    // rom_array[21652] = 32'hFFFFFFF0;
    // rom_array[21653] = 32'hFFFFFFF1;
    // rom_array[21654] = 32'hFFFFFFF1;
    // rom_array[21655] = 32'hFFFFFFF1;
    // rom_array[21656] = 32'hFFFFFFF1;
    // rom_array[21657] = 32'hFFFFFFF1;
    // rom_array[21658] = 32'hFFFFFFF1;
    // rom_array[21659] = 32'hFFFFFFF1;
    // rom_array[21660] = 32'hFFFFFFF1;
    // rom_array[21661] = 32'hFFFFFFF1;
    // rom_array[21662] = 32'hFFFFFFF1;
    // rom_array[21663] = 32'hFFFFFFF1;
    // rom_array[21664] = 32'hFFFFFFF1;
    // rom_array[21665] = 32'hFFFFFFF1;
    // rom_array[21666] = 32'hFFFFFFF1;
    // rom_array[21667] = 32'hFFFFFFF1;
    // rom_array[21668] = 32'hFFFFFFF1;
    // rom_array[21669] = 32'hFFFFFFF1;
    // rom_array[21670] = 32'hFFFFFFF1;
    // rom_array[21671] = 32'hFFFFFFF1;
    // rom_array[21672] = 32'hFFFFFFF1;
    // rom_array[21673] = 32'hFFFFFFF1;
    // rom_array[21674] = 32'hFFFFFFF1;
    // rom_array[21675] = 32'hFFFFFFF1;
    // rom_array[21676] = 32'hFFFFFFF1;
    // rom_array[21677] = 32'hFFFFFFF1;
    // rom_array[21678] = 32'hFFFFFFF1;
    // rom_array[21679] = 32'hFFFFFFF1;
    // rom_array[21680] = 32'hFFFFFFF1;
    // rom_array[21681] = 32'hFFFFFFF1;
    // rom_array[21682] = 32'hFFFFFFF1;
    // rom_array[21683] = 32'hFFFFFFF1;
    // rom_array[21684] = 32'hFFFFFFF1;
    // rom_array[21685] = 32'hFFFFFFF1;
    // rom_array[21686] = 32'hFFFFFFF1;
    // rom_array[21687] = 32'hFFFFFFF1;
    // rom_array[21688] = 32'hFFFFFFF1;
    // rom_array[21689] = 32'hFFFFFFF0;
    // rom_array[21690] = 32'hFFFFFFF0;
    // rom_array[21691] = 32'hFFFFFFF0;
    // rom_array[21692] = 32'hFFFFFFF0;
    // rom_array[21693] = 32'hFFFFFFF1;
    // rom_array[21694] = 32'hFFFFFFF1;
    // rom_array[21695] = 32'hFFFFFFF1;
    // rom_array[21696] = 32'hFFFFFFF1;
    // rom_array[21697] = 32'hFFFFFFF0;
    // rom_array[21698] = 32'hFFFFFFF0;
    // rom_array[21699] = 32'hFFFFFFF0;
    // rom_array[21700] = 32'hFFFFFFF0;
    // rom_array[21701] = 32'hFFFFFFF1;
    // rom_array[21702] = 32'hFFFFFFF1;
    // rom_array[21703] = 32'hFFFFFFF1;
    // rom_array[21704] = 32'hFFFFFFF1;
    // rom_array[21705] = 32'hFFFFFFF0;
    // rom_array[21706] = 32'hFFFFFFF0;
    // rom_array[21707] = 32'hFFFFFFF0;
    // rom_array[21708] = 32'hFFFFFFF0;
    // rom_array[21709] = 32'hFFFFFFF1;
    // rom_array[21710] = 32'hFFFFFFF1;
    // rom_array[21711] = 32'hFFFFFFF1;
    // rom_array[21712] = 32'hFFFFFFF1;
    // rom_array[21713] = 32'hFFFFFFF0;
    // rom_array[21714] = 32'hFFFFFFF0;
    // rom_array[21715] = 32'hFFFFFFF0;
    // rom_array[21716] = 32'hFFFFFFF0;
    // rom_array[21717] = 32'hFFFFFFF1;
    // rom_array[21718] = 32'hFFFFFFF1;
    // rom_array[21719] = 32'hFFFFFFF1;
    // rom_array[21720] = 32'hFFFFFFF1;
    // rom_array[21721] = 32'hFFFFFFF1;
    // rom_array[21722] = 32'hFFFFFFF1;
    // rom_array[21723] = 32'hFFFFFFF1;
    // rom_array[21724] = 32'hFFFFFFF1;
    // rom_array[21725] = 32'hFFFFFFF1;
    // rom_array[21726] = 32'hFFFFFFF1;
    // rom_array[21727] = 32'hFFFFFFF1;
    // rom_array[21728] = 32'hFFFFFFF1;
    // rom_array[21729] = 32'hFFFFFFF1;
    // rom_array[21730] = 32'hFFFFFFF1;
    // rom_array[21731] = 32'hFFFFFFF1;
    // rom_array[21732] = 32'hFFFFFFF1;
    // rom_array[21733] = 32'hFFFFFFF1;
    // rom_array[21734] = 32'hFFFFFFF1;
    // rom_array[21735] = 32'hFFFFFFF1;
    // rom_array[21736] = 32'hFFFFFFF1;
    // rom_array[21737] = 32'hFFFFFFF1;
    // rom_array[21738] = 32'hFFFFFFF1;
    // rom_array[21739] = 32'hFFFFFFF1;
    // rom_array[21740] = 32'hFFFFFFF1;
    // rom_array[21741] = 32'hFFFFFFF1;
    // rom_array[21742] = 32'hFFFFFFF1;
    // rom_array[21743] = 32'hFFFFFFF1;
    // rom_array[21744] = 32'hFFFFFFF1;
    // rom_array[21745] = 32'hFFFFFFF1;
    // rom_array[21746] = 32'hFFFFFFF1;
    // rom_array[21747] = 32'hFFFFFFF1;
    // rom_array[21748] = 32'hFFFFFFF1;
    // rom_array[21749] = 32'hFFFFFFF1;
    // rom_array[21750] = 32'hFFFFFFF1;
    // rom_array[21751] = 32'hFFFFFFF1;
    // rom_array[21752] = 32'hFFFFFFF1;
    // rom_array[21753] = 32'hFFFFFFF0;
    // rom_array[21754] = 32'hFFFFFFF0;
    // rom_array[21755] = 32'hFFFFFFF0;
    // rom_array[21756] = 32'hFFFFFFF0;
    // rom_array[21757] = 32'hFFFFFFF1;
    // rom_array[21758] = 32'hFFFFFFF1;
    // rom_array[21759] = 32'hFFFFFFF1;
    // rom_array[21760] = 32'hFFFFFFF1;
    // rom_array[21761] = 32'hFFFFFFF0;
    // rom_array[21762] = 32'hFFFFFFF0;
    // rom_array[21763] = 32'hFFFFFFF0;
    // rom_array[21764] = 32'hFFFFFFF0;
    // rom_array[21765] = 32'hFFFFFFF1;
    // rom_array[21766] = 32'hFFFFFFF1;
    // rom_array[21767] = 32'hFFFFFFF1;
    // rom_array[21768] = 32'hFFFFFFF1;
    // rom_array[21769] = 32'hFFFFFFF0;
    // rom_array[21770] = 32'hFFFFFFF0;
    // rom_array[21771] = 32'hFFFFFFF0;
    // rom_array[21772] = 32'hFFFFFFF0;
    // rom_array[21773] = 32'hFFFFFFF1;
    // rom_array[21774] = 32'hFFFFFFF1;
    // rom_array[21775] = 32'hFFFFFFF1;
    // rom_array[21776] = 32'hFFFFFFF1;
    // rom_array[21777] = 32'hFFFFFFF0;
    // rom_array[21778] = 32'hFFFFFFF0;
    // rom_array[21779] = 32'hFFFFFFF0;
    // rom_array[21780] = 32'hFFFFFFF0;
    // rom_array[21781] = 32'hFFFFFFF1;
    // rom_array[21782] = 32'hFFFFFFF1;
    // rom_array[21783] = 32'hFFFFFFF1;
    // rom_array[21784] = 32'hFFFFFFF1;
    // rom_array[21785] = 32'hFFFFFFF1;
    // rom_array[21786] = 32'hFFFFFFF1;
    // rom_array[21787] = 32'hFFFFFFF1;
    // rom_array[21788] = 32'hFFFFFFF1;
    // rom_array[21789] = 32'hFFFFFFF1;
    // rom_array[21790] = 32'hFFFFFFF1;
    // rom_array[21791] = 32'hFFFFFFF1;
    // rom_array[21792] = 32'hFFFFFFF1;
    // rom_array[21793] = 32'hFFFFFFF1;
    // rom_array[21794] = 32'hFFFFFFF1;
    // rom_array[21795] = 32'hFFFFFFF1;
    // rom_array[21796] = 32'hFFFFFFF1;
    // rom_array[21797] = 32'hFFFFFFF1;
    // rom_array[21798] = 32'hFFFFFFF1;
    // rom_array[21799] = 32'hFFFFFFF1;
    // rom_array[21800] = 32'hFFFFFFF1;
    // rom_array[21801] = 32'hFFFFFFF1;
    // rom_array[21802] = 32'hFFFFFFF1;
    // rom_array[21803] = 32'hFFFFFFF1;
    // rom_array[21804] = 32'hFFFFFFF1;
    // rom_array[21805] = 32'hFFFFFFF1;
    // rom_array[21806] = 32'hFFFFFFF1;
    // rom_array[21807] = 32'hFFFFFFF1;
    // rom_array[21808] = 32'hFFFFFFF1;
    // rom_array[21809] = 32'hFFFFFFF1;
    // rom_array[21810] = 32'hFFFFFFF1;
    // rom_array[21811] = 32'hFFFFFFF1;
    // rom_array[21812] = 32'hFFFFFFF1;
    // rom_array[21813] = 32'hFFFFFFF1;
    // rom_array[21814] = 32'hFFFFFFF1;
    // rom_array[21815] = 32'hFFFFFFF1;
    // rom_array[21816] = 32'hFFFFFFF1;
    // rom_array[21817] = 32'hFFFFFFF0;
    // rom_array[21818] = 32'hFFFFFFF0;
    // rom_array[21819] = 32'hFFFFFFF0;
    // rom_array[21820] = 32'hFFFFFFF0;
    // rom_array[21821] = 32'hFFFFFFF1;
    // rom_array[21822] = 32'hFFFFFFF1;
    // rom_array[21823] = 32'hFFFFFFF1;
    // rom_array[21824] = 32'hFFFFFFF1;
    // rom_array[21825] = 32'hFFFFFFF0;
    // rom_array[21826] = 32'hFFFFFFF0;
    // rom_array[21827] = 32'hFFFFFFF0;
    // rom_array[21828] = 32'hFFFFFFF0;
    // rom_array[21829] = 32'hFFFFFFF1;
    // rom_array[21830] = 32'hFFFFFFF1;
    // rom_array[21831] = 32'hFFFFFFF1;
    // rom_array[21832] = 32'hFFFFFFF1;
    // rom_array[21833] = 32'hFFFFFFF0;
    // rom_array[21834] = 32'hFFFFFFF0;
    // rom_array[21835] = 32'hFFFFFFF0;
    // rom_array[21836] = 32'hFFFFFFF0;
    // rom_array[21837] = 32'hFFFFFFF1;
    // rom_array[21838] = 32'hFFFFFFF1;
    // rom_array[21839] = 32'hFFFFFFF1;
    // rom_array[21840] = 32'hFFFFFFF1;
    // rom_array[21841] = 32'hFFFFFFF0;
    // rom_array[21842] = 32'hFFFFFFF0;
    // rom_array[21843] = 32'hFFFFFFF0;
    // rom_array[21844] = 32'hFFFFFFF0;
    // rom_array[21845] = 32'hFFFFFFF1;
    // rom_array[21846] = 32'hFFFFFFF1;
    // rom_array[21847] = 32'hFFFFFFF1;
    // rom_array[21848] = 32'hFFFFFFF1;
    // rom_array[21849] = 32'hFFFFFFF1;
    // rom_array[21850] = 32'hFFFFFFF1;
    // rom_array[21851] = 32'hFFFFFFF1;
    // rom_array[21852] = 32'hFFFFFFF1;
    // rom_array[21853] = 32'hFFFFFFF1;
    // rom_array[21854] = 32'hFFFFFFF1;
    // rom_array[21855] = 32'hFFFFFFF1;
    // rom_array[21856] = 32'hFFFFFFF1;
    // rom_array[21857] = 32'hFFFFFFF1;
    // rom_array[21858] = 32'hFFFFFFF1;
    // rom_array[21859] = 32'hFFFFFFF1;
    // rom_array[21860] = 32'hFFFFFFF1;
    // rom_array[21861] = 32'hFFFFFFF1;
    // rom_array[21862] = 32'hFFFFFFF1;
    // rom_array[21863] = 32'hFFFFFFF1;
    // rom_array[21864] = 32'hFFFFFFF1;
    // rom_array[21865] = 32'hFFFFFFF1;
    // rom_array[21866] = 32'hFFFFFFF1;
    // rom_array[21867] = 32'hFFFFFFF1;
    // rom_array[21868] = 32'hFFFFFFF1;
    // rom_array[21869] = 32'hFFFFFFF1;
    // rom_array[21870] = 32'hFFFFFFF1;
    // rom_array[21871] = 32'hFFFFFFF1;
    // rom_array[21872] = 32'hFFFFFFF1;
    // rom_array[21873] = 32'hFFFFFFF1;
    // rom_array[21874] = 32'hFFFFFFF1;
    // rom_array[21875] = 32'hFFFFFFF1;
    // rom_array[21876] = 32'hFFFFFFF1;
    // rom_array[21877] = 32'hFFFFFFF1;
    // rom_array[21878] = 32'hFFFFFFF1;
    // rom_array[21879] = 32'hFFFFFFF1;
    // rom_array[21880] = 32'hFFFFFFF1;
    // rom_array[21881] = 32'hFFFFFFF0;
    // rom_array[21882] = 32'hFFFFFFF0;
    // rom_array[21883] = 32'hFFFFFFF0;
    // rom_array[21884] = 32'hFFFFFFF0;
    // rom_array[21885] = 32'hFFFFFFF1;
    // rom_array[21886] = 32'hFFFFFFF1;
    // rom_array[21887] = 32'hFFFFFFF1;
    // rom_array[21888] = 32'hFFFFFFF1;
    // rom_array[21889] = 32'hFFFFFFF0;
    // rom_array[21890] = 32'hFFFFFFF0;
    // rom_array[21891] = 32'hFFFFFFF0;
    // rom_array[21892] = 32'hFFFFFFF0;
    // rom_array[21893] = 32'hFFFFFFF1;
    // rom_array[21894] = 32'hFFFFFFF1;
    // rom_array[21895] = 32'hFFFFFFF1;
    // rom_array[21896] = 32'hFFFFFFF1;
    // rom_array[21897] = 32'hFFFFFFF0;
    // rom_array[21898] = 32'hFFFFFFF0;
    // rom_array[21899] = 32'hFFFFFFF0;
    // rom_array[21900] = 32'hFFFFFFF0;
    // rom_array[21901] = 32'hFFFFFFF1;
    // rom_array[21902] = 32'hFFFFFFF1;
    // rom_array[21903] = 32'hFFFFFFF1;
    // rom_array[21904] = 32'hFFFFFFF1;
    // rom_array[21905] = 32'hFFFFFFF0;
    // rom_array[21906] = 32'hFFFFFFF0;
    // rom_array[21907] = 32'hFFFFFFF0;
    // rom_array[21908] = 32'hFFFFFFF0;
    // rom_array[21909] = 32'hFFFFFFF1;
    // rom_array[21910] = 32'hFFFFFFF1;
    // rom_array[21911] = 32'hFFFFFFF1;
    // rom_array[21912] = 32'hFFFFFFF1;
    // rom_array[21913] = 32'hFFFFFFF1;
    // rom_array[21914] = 32'hFFFFFFF1;
    // rom_array[21915] = 32'hFFFFFFF1;
    // rom_array[21916] = 32'hFFFFFFF1;
    // rom_array[21917] = 32'hFFFFFFF1;
    // rom_array[21918] = 32'hFFFFFFF1;
    // rom_array[21919] = 32'hFFFFFFF1;
    // rom_array[21920] = 32'hFFFFFFF1;
    // rom_array[21921] = 32'hFFFFFFF1;
    // rom_array[21922] = 32'hFFFFFFF1;
    // rom_array[21923] = 32'hFFFFFFF1;
    // rom_array[21924] = 32'hFFFFFFF1;
    // rom_array[21925] = 32'hFFFFFFF1;
    // rom_array[21926] = 32'hFFFFFFF1;
    // rom_array[21927] = 32'hFFFFFFF1;
    // rom_array[21928] = 32'hFFFFFFF1;
    // rom_array[21929] = 32'hFFFFFFF1;
    // rom_array[21930] = 32'hFFFFFFF1;
    // rom_array[21931] = 32'hFFFFFFF1;
    // rom_array[21932] = 32'hFFFFFFF1;
    // rom_array[21933] = 32'hFFFFFFF1;
    // rom_array[21934] = 32'hFFFFFFF1;
    // rom_array[21935] = 32'hFFFFFFF1;
    // rom_array[21936] = 32'hFFFFFFF1;
    // rom_array[21937] = 32'hFFFFFFF1;
    // rom_array[21938] = 32'hFFFFFFF1;
    // rom_array[21939] = 32'hFFFFFFF1;
    // rom_array[21940] = 32'hFFFFFFF1;
    // rom_array[21941] = 32'hFFFFFFF1;
    // rom_array[21942] = 32'hFFFFFFF1;
    // rom_array[21943] = 32'hFFFFFFF1;
    // rom_array[21944] = 32'hFFFFFFF1;
    // rom_array[21945] = 32'hFFFFFFF0;
    // rom_array[21946] = 32'hFFFFFFF0;
    // rom_array[21947] = 32'hFFFFFFF0;
    // rom_array[21948] = 32'hFFFFFFF0;
    // rom_array[21949] = 32'hFFFFFFF1;
    // rom_array[21950] = 32'hFFFFFFF1;
    // rom_array[21951] = 32'hFFFFFFF1;
    // rom_array[21952] = 32'hFFFFFFF1;
    // rom_array[21953] = 32'hFFFFFFF0;
    // rom_array[21954] = 32'hFFFFFFF0;
    // rom_array[21955] = 32'hFFFFFFF0;
    // rom_array[21956] = 32'hFFFFFFF0;
    // rom_array[21957] = 32'hFFFFFFF1;
    // rom_array[21958] = 32'hFFFFFFF1;
    // rom_array[21959] = 32'hFFFFFFF1;
    // rom_array[21960] = 32'hFFFFFFF1;
    // rom_array[21961] = 32'hFFFFFFF1;
    // rom_array[21962] = 32'hFFFFFFF1;
    // rom_array[21963] = 32'hFFFFFFF1;
    // rom_array[21964] = 32'hFFFFFFF1;
    // rom_array[21965] = 32'hFFFFFFF1;
    // rom_array[21966] = 32'hFFFFFFF1;
    // rom_array[21967] = 32'hFFFFFFF1;
    // rom_array[21968] = 32'hFFFFFFF1;
    // rom_array[21969] = 32'hFFFFFFF1;
    // rom_array[21970] = 32'hFFFFFFF1;
    // rom_array[21971] = 32'hFFFFFFF1;
    // rom_array[21972] = 32'hFFFFFFF1;
    // rom_array[21973] = 32'hFFFFFFF1;
    // rom_array[21974] = 32'hFFFFFFF1;
    // rom_array[21975] = 32'hFFFFFFF1;
    // rom_array[21976] = 32'hFFFFFFF1;
    // rom_array[21977] = 32'hFFFFFFF1;
    // rom_array[21978] = 32'hFFFFFFF1;
    // rom_array[21979] = 32'hFFFFFFF0;
    // rom_array[21980] = 32'hFFFFFFF0;
    // rom_array[21981] = 32'hFFFFFFF1;
    // rom_array[21982] = 32'hFFFFFFF1;
    // rom_array[21983] = 32'hFFFFFFF0;
    // rom_array[21984] = 32'hFFFFFFF0;
    // rom_array[21985] = 32'hFFFFFFF1;
    // rom_array[21986] = 32'hFFFFFFF1;
    // rom_array[21987] = 32'hFFFFFFF0;
    // rom_array[21988] = 32'hFFFFFFF0;
    // rom_array[21989] = 32'hFFFFFFF1;
    // rom_array[21990] = 32'hFFFFFFF1;
    // rom_array[21991] = 32'hFFFFFFF0;
    // rom_array[21992] = 32'hFFFFFFF0;
    // rom_array[21993] = 32'hFFFFFFF1;
    // rom_array[21994] = 32'hFFFFFFF1;
    // rom_array[21995] = 32'hFFFFFFF1;
    // rom_array[21996] = 32'hFFFFFFF1;
    // rom_array[21997] = 32'hFFFFFFF0;
    // rom_array[21998] = 32'hFFFFFFF0;
    // rom_array[21999] = 32'hFFFFFFF0;
    // rom_array[22000] = 32'hFFFFFFF0;
    // rom_array[22001] = 32'hFFFFFFF1;
    // rom_array[22002] = 32'hFFFFFFF1;
    // rom_array[22003] = 32'hFFFFFFF1;
    // rom_array[22004] = 32'hFFFFFFF1;
    // rom_array[22005] = 32'hFFFFFFF0;
    // rom_array[22006] = 32'hFFFFFFF0;
    // rom_array[22007] = 32'hFFFFFFF0;
    // rom_array[22008] = 32'hFFFFFFF0;
    // rom_array[22009] = 32'hFFFFFFF1;
    // rom_array[22010] = 32'hFFFFFFF1;
    // rom_array[22011] = 32'hFFFFFFF1;
    // rom_array[22012] = 32'hFFFFFFF1;
    // rom_array[22013] = 32'hFFFFFFF0;
    // rom_array[22014] = 32'hFFFFFFF0;
    // rom_array[22015] = 32'hFFFFFFF0;
    // rom_array[22016] = 32'hFFFFFFF0;
    // rom_array[22017] = 32'hFFFFFFF1;
    // rom_array[22018] = 32'hFFFFFFF1;
    // rom_array[22019] = 32'hFFFFFFF1;
    // rom_array[22020] = 32'hFFFFFFF1;
    // rom_array[22021] = 32'hFFFFFFF0;
    // rom_array[22022] = 32'hFFFFFFF0;
    // rom_array[22023] = 32'hFFFFFFF0;
    // rom_array[22024] = 32'hFFFFFFF0;
    // rom_array[22025] = 32'hFFFFFFF1;
    // rom_array[22026] = 32'hFFFFFFF1;
    // rom_array[22027] = 32'hFFFFFFF1;
    // rom_array[22028] = 32'hFFFFFFF1;
    // rom_array[22029] = 32'hFFFFFFF0;
    // rom_array[22030] = 32'hFFFFFFF0;
    // rom_array[22031] = 32'hFFFFFFF0;
    // rom_array[22032] = 32'hFFFFFFF0;
    // rom_array[22033] = 32'hFFFFFFF1;
    // rom_array[22034] = 32'hFFFFFFF1;
    // rom_array[22035] = 32'hFFFFFFF1;
    // rom_array[22036] = 32'hFFFFFFF1;
    // rom_array[22037] = 32'hFFFFFFF0;
    // rom_array[22038] = 32'hFFFFFFF0;
    // rom_array[22039] = 32'hFFFFFFF0;
    // rom_array[22040] = 32'hFFFFFFF0;
    // rom_array[22041] = 32'hFFFFFFF1;
    // rom_array[22042] = 32'hFFFFFFF1;
    // rom_array[22043] = 32'hFFFFFFF1;
    // rom_array[22044] = 32'hFFFFFFF1;
    // rom_array[22045] = 32'hFFFFFFF0;
    // rom_array[22046] = 32'hFFFFFFF0;
    // rom_array[22047] = 32'hFFFFFFF0;
    // rom_array[22048] = 32'hFFFFFFF0;
    // rom_array[22049] = 32'hFFFFFFF1;
    // rom_array[22050] = 32'hFFFFFFF1;
    // rom_array[22051] = 32'hFFFFFFF1;
    // rom_array[22052] = 32'hFFFFFFF1;
    // rom_array[22053] = 32'hFFFFFFF0;
    // rom_array[22054] = 32'hFFFFFFF0;
    // rom_array[22055] = 32'hFFFFFFF0;
    // rom_array[22056] = 32'hFFFFFFF0;
    // rom_array[22057] = 32'hFFFFFFF1;
    // rom_array[22058] = 32'hFFFFFFF1;
    // rom_array[22059] = 32'hFFFFFFF1;
    // rom_array[22060] = 32'hFFFFFFF1;
    // rom_array[22061] = 32'hFFFFFFF0;
    // rom_array[22062] = 32'hFFFFFFF0;
    // rom_array[22063] = 32'hFFFFFFF0;
    // rom_array[22064] = 32'hFFFFFFF0;
    // rom_array[22065] = 32'hFFFFFFF1;
    // rom_array[22066] = 32'hFFFFFFF1;
    // rom_array[22067] = 32'hFFFFFFF1;
    // rom_array[22068] = 32'hFFFFFFF1;
    // rom_array[22069] = 32'hFFFFFFF0;
    // rom_array[22070] = 32'hFFFFFFF0;
    // rom_array[22071] = 32'hFFFFFFF0;
    // rom_array[22072] = 32'hFFFFFFF0;
    // rom_array[22073] = 32'hFFFFFFF1;
    // rom_array[22074] = 32'hFFFFFFF1;
    // rom_array[22075] = 32'hFFFFFFF1;
    // rom_array[22076] = 32'hFFFFFFF1;
    // rom_array[22077] = 32'hFFFFFFF0;
    // rom_array[22078] = 32'hFFFFFFF0;
    // rom_array[22079] = 32'hFFFFFFF0;
    // rom_array[22080] = 32'hFFFFFFF0;
    // rom_array[22081] = 32'hFFFFFFF1;
    // rom_array[22082] = 32'hFFFFFFF1;
    // rom_array[22083] = 32'hFFFFFFF1;
    // rom_array[22084] = 32'hFFFFFFF1;
    // rom_array[22085] = 32'hFFFFFFF0;
    // rom_array[22086] = 32'hFFFFFFF0;
    // rom_array[22087] = 32'hFFFFFFF0;
    // rom_array[22088] = 32'hFFFFFFF0;
    // rom_array[22089] = 32'hFFFFFFF1;
    // rom_array[22090] = 32'hFFFFFFF1;
    // rom_array[22091] = 32'hFFFFFFF1;
    // rom_array[22092] = 32'hFFFFFFF1;
    // rom_array[22093] = 32'hFFFFFFF0;
    // rom_array[22094] = 32'hFFFFFFF0;
    // rom_array[22095] = 32'hFFFFFFF0;
    // rom_array[22096] = 32'hFFFFFFF0;
    // rom_array[22097] = 32'hFFFFFFF1;
    // rom_array[22098] = 32'hFFFFFFF1;
    // rom_array[22099] = 32'hFFFFFFF1;
    // rom_array[22100] = 32'hFFFFFFF1;
    // rom_array[22101] = 32'hFFFFFFF0;
    // rom_array[22102] = 32'hFFFFFFF0;
    // rom_array[22103] = 32'hFFFFFFF0;
    // rom_array[22104] = 32'hFFFFFFF0;
    // rom_array[22105] = 32'hFFFFFFF1;
    // rom_array[22106] = 32'hFFFFFFF1;
    // rom_array[22107] = 32'hFFFFFFF1;
    // rom_array[22108] = 32'hFFFFFFF1;
    // rom_array[22109] = 32'hFFFFFFF0;
    // rom_array[22110] = 32'hFFFFFFF0;
    // rom_array[22111] = 32'hFFFFFFF0;
    // rom_array[22112] = 32'hFFFFFFF0;
    // rom_array[22113] = 32'hFFFFFFF1;
    // rom_array[22114] = 32'hFFFFFFF1;
    // rom_array[22115] = 32'hFFFFFFF1;
    // rom_array[22116] = 32'hFFFFFFF1;
    // rom_array[22117] = 32'hFFFFFFF0;
    // rom_array[22118] = 32'hFFFFFFF0;
    // rom_array[22119] = 32'hFFFFFFF0;
    // rom_array[22120] = 32'hFFFFFFF0;
    // rom_array[22121] = 32'hFFFFFFF1;
    // rom_array[22122] = 32'hFFFFFFF1;
    // rom_array[22123] = 32'hFFFFFFF1;
    // rom_array[22124] = 32'hFFFFFFF1;
    // rom_array[22125] = 32'hFFFFFFF1;
    // rom_array[22126] = 32'hFFFFFFF1;
    // rom_array[22127] = 32'hFFFFFFF1;
    // rom_array[22128] = 32'hFFFFFFF1;
    // rom_array[22129] = 32'hFFFFFFF1;
    // rom_array[22130] = 32'hFFFFFFF1;
    // rom_array[22131] = 32'hFFFFFFF1;
    // rom_array[22132] = 32'hFFFFFFF1;
    // rom_array[22133] = 32'hFFFFFFF1;
    // rom_array[22134] = 32'hFFFFFFF1;
    // rom_array[22135] = 32'hFFFFFFF1;
    // rom_array[22136] = 32'hFFFFFFF1;
    // rom_array[22137] = 32'hFFFFFFF1;
    // rom_array[22138] = 32'hFFFFFFF1;
    // rom_array[22139] = 32'hFFFFFFF0;
    // rom_array[22140] = 32'hFFFFFFF0;
    // rom_array[22141] = 32'hFFFFFFF1;
    // rom_array[22142] = 32'hFFFFFFF1;
    // rom_array[22143] = 32'hFFFFFFF0;
    // rom_array[22144] = 32'hFFFFFFF0;
    // rom_array[22145] = 32'hFFFFFFF1;
    // rom_array[22146] = 32'hFFFFFFF1;
    // rom_array[22147] = 32'hFFFFFFF0;
    // rom_array[22148] = 32'hFFFFFFF0;
    // rom_array[22149] = 32'hFFFFFFF1;
    // rom_array[22150] = 32'hFFFFFFF1;
    // rom_array[22151] = 32'hFFFFFFF0;
    // rom_array[22152] = 32'hFFFFFFF0;
    // rom_array[22153] = 32'hFFFFFFF1;
    // rom_array[22154] = 32'hFFFFFFF1;
    // rom_array[22155] = 32'hFFFFFFF1;
    // rom_array[22156] = 32'hFFFFFFF1;
    // rom_array[22157] = 32'hFFFFFFF1;
    // rom_array[22158] = 32'hFFFFFFF1;
    // rom_array[22159] = 32'hFFFFFFF1;
    // rom_array[22160] = 32'hFFFFFFF1;
    // rom_array[22161] = 32'hFFFFFFF1;
    // rom_array[22162] = 32'hFFFFFFF1;
    // rom_array[22163] = 32'hFFFFFFF1;
    // rom_array[22164] = 32'hFFFFFFF1;
    // rom_array[22165] = 32'hFFFFFFF1;
    // rom_array[22166] = 32'hFFFFFFF1;
    // rom_array[22167] = 32'hFFFFFFF1;
    // rom_array[22168] = 32'hFFFFFFF1;
    // rom_array[22169] = 32'hFFFFFFF1;
    // rom_array[22170] = 32'hFFFFFFF1;
    // rom_array[22171] = 32'hFFFFFFF0;
    // rom_array[22172] = 32'hFFFFFFF0;
    // rom_array[22173] = 32'hFFFFFFF1;
    // rom_array[22174] = 32'hFFFFFFF1;
    // rom_array[22175] = 32'hFFFFFFF0;
    // rom_array[22176] = 32'hFFFFFFF0;
    // rom_array[22177] = 32'hFFFFFFF1;
    // rom_array[22178] = 32'hFFFFFFF1;
    // rom_array[22179] = 32'hFFFFFFF0;
    // rom_array[22180] = 32'hFFFFFFF0;
    // rom_array[22181] = 32'hFFFFFFF1;
    // rom_array[22182] = 32'hFFFFFFF1;
    // rom_array[22183] = 32'hFFFFFFF0;
    // rom_array[22184] = 32'hFFFFFFF0;
    // rom_array[22185] = 32'hFFFFFFF1;
    // rom_array[22186] = 32'hFFFFFFF1;
    // rom_array[22187] = 32'hFFFFFFF1;
    // rom_array[22188] = 32'hFFFFFFF1;
    // rom_array[22189] = 32'hFFFFFFF0;
    // rom_array[22190] = 32'hFFFFFFF0;
    // rom_array[22191] = 32'hFFFFFFF0;
    // rom_array[22192] = 32'hFFFFFFF0;
    // rom_array[22193] = 32'hFFFFFFF1;
    // rom_array[22194] = 32'hFFFFFFF1;
    // rom_array[22195] = 32'hFFFFFFF1;
    // rom_array[22196] = 32'hFFFFFFF1;
    // rom_array[22197] = 32'hFFFFFFF0;
    // rom_array[22198] = 32'hFFFFFFF0;
    // rom_array[22199] = 32'hFFFFFFF0;
    // rom_array[22200] = 32'hFFFFFFF0;
    // rom_array[22201] = 32'hFFFFFFF1;
    // rom_array[22202] = 32'hFFFFFFF1;
    // rom_array[22203] = 32'hFFFFFFF1;
    // rom_array[22204] = 32'hFFFFFFF1;
    // rom_array[22205] = 32'hFFFFFFF0;
    // rom_array[22206] = 32'hFFFFFFF0;
    // rom_array[22207] = 32'hFFFFFFF0;
    // rom_array[22208] = 32'hFFFFFFF0;
    // rom_array[22209] = 32'hFFFFFFF1;
    // rom_array[22210] = 32'hFFFFFFF1;
    // rom_array[22211] = 32'hFFFFFFF1;
    // rom_array[22212] = 32'hFFFFFFF1;
    // rom_array[22213] = 32'hFFFFFFF0;
    // rom_array[22214] = 32'hFFFFFFF0;
    // rom_array[22215] = 32'hFFFFFFF0;
    // rom_array[22216] = 32'hFFFFFFF0;
    // rom_array[22217] = 32'hFFFFFFF1;
    // rom_array[22218] = 32'hFFFFFFF1;
    // rom_array[22219] = 32'hFFFFFFF1;
    // rom_array[22220] = 32'hFFFFFFF1;
    // rom_array[22221] = 32'hFFFFFFF0;
    // rom_array[22222] = 32'hFFFFFFF0;
    // rom_array[22223] = 32'hFFFFFFF0;
    // rom_array[22224] = 32'hFFFFFFF0;
    // rom_array[22225] = 32'hFFFFFFF1;
    // rom_array[22226] = 32'hFFFFFFF1;
    // rom_array[22227] = 32'hFFFFFFF1;
    // rom_array[22228] = 32'hFFFFFFF1;
    // rom_array[22229] = 32'hFFFFFFF0;
    // rom_array[22230] = 32'hFFFFFFF0;
    // rom_array[22231] = 32'hFFFFFFF0;
    // rom_array[22232] = 32'hFFFFFFF0;
    // rom_array[22233] = 32'hFFFFFFF1;
    // rom_array[22234] = 32'hFFFFFFF1;
    // rom_array[22235] = 32'hFFFFFFF0;
    // rom_array[22236] = 32'hFFFFFFF0;
    // rom_array[22237] = 32'hFFFFFFF1;
    // rom_array[22238] = 32'hFFFFFFF1;
    // rom_array[22239] = 32'hFFFFFFF0;
    // rom_array[22240] = 32'hFFFFFFF0;
    // rom_array[22241] = 32'hFFFFFFF1;
    // rom_array[22242] = 32'hFFFFFFF1;
    // rom_array[22243] = 32'hFFFFFFF0;
    // rom_array[22244] = 32'hFFFFFFF0;
    // rom_array[22245] = 32'hFFFFFFF1;
    // rom_array[22246] = 32'hFFFFFFF1;
    // rom_array[22247] = 32'hFFFFFFF0;
    // rom_array[22248] = 32'hFFFFFFF0;
    // rom_array[22249] = 32'hFFFFFFF1;
    // rom_array[22250] = 32'hFFFFFFF1;
    // rom_array[22251] = 32'hFFFFFFF0;
    // rom_array[22252] = 32'hFFFFFFF0;
    // rom_array[22253] = 32'hFFFFFFF1;
    // rom_array[22254] = 32'hFFFFFFF1;
    // rom_array[22255] = 32'hFFFFFFF0;
    // rom_array[22256] = 32'hFFFFFFF0;
    // rom_array[22257] = 32'hFFFFFFF1;
    // rom_array[22258] = 32'hFFFFFFF1;
    // rom_array[22259] = 32'hFFFFFFF0;
    // rom_array[22260] = 32'hFFFFFFF0;
    // rom_array[22261] = 32'hFFFFFFF1;
    // rom_array[22262] = 32'hFFFFFFF1;
    // rom_array[22263] = 32'hFFFFFFF0;
    // rom_array[22264] = 32'hFFFFFFF0;
    // rom_array[22265] = 32'hFFFFFFF1;
    // rom_array[22266] = 32'hFFFFFFF1;
    // rom_array[22267] = 32'hFFFFFFF0;
    // rom_array[22268] = 32'hFFFFFFF0;
    // rom_array[22269] = 32'hFFFFFFF1;
    // rom_array[22270] = 32'hFFFFFFF1;
    // rom_array[22271] = 32'hFFFFFFF0;
    // rom_array[22272] = 32'hFFFFFFF0;
    // rom_array[22273] = 32'hFFFFFFF1;
    // rom_array[22274] = 32'hFFFFFFF1;
    // rom_array[22275] = 32'hFFFFFFF0;
    // rom_array[22276] = 32'hFFFFFFF0;
    // rom_array[22277] = 32'hFFFFFFF1;
    // rom_array[22278] = 32'hFFFFFFF1;
    // rom_array[22279] = 32'hFFFFFFF0;
    // rom_array[22280] = 32'hFFFFFFF0;
    // rom_array[22281] = 32'hFFFFFFF1;
    // rom_array[22282] = 32'hFFFFFFF1;
    // rom_array[22283] = 32'hFFFFFFF0;
    // rom_array[22284] = 32'hFFFFFFF0;
    // rom_array[22285] = 32'hFFFFFFF1;
    // rom_array[22286] = 32'hFFFFFFF1;
    // rom_array[22287] = 32'hFFFFFFF0;
    // rom_array[22288] = 32'hFFFFFFF0;
    // rom_array[22289] = 32'hFFFFFFF1;
    // rom_array[22290] = 32'hFFFFFFF1;
    // rom_array[22291] = 32'hFFFFFFF0;
    // rom_array[22292] = 32'hFFFFFFF0;
    // rom_array[22293] = 32'hFFFFFFF1;
    // rom_array[22294] = 32'hFFFFFFF1;
    // rom_array[22295] = 32'hFFFFFFF0;
    // rom_array[22296] = 32'hFFFFFFF0;
    // rom_array[22297] = 32'hFFFFFFF1;
    // rom_array[22298] = 32'hFFFFFFF1;
    // rom_array[22299] = 32'hFFFFFFF0;
    // rom_array[22300] = 32'hFFFFFFF0;
    // rom_array[22301] = 32'hFFFFFFF1;
    // rom_array[22302] = 32'hFFFFFFF1;
    // rom_array[22303] = 32'hFFFFFFF0;
    // rom_array[22304] = 32'hFFFFFFF0;
    // rom_array[22305] = 32'hFFFFFFF1;
    // rom_array[22306] = 32'hFFFFFFF1;
    // rom_array[22307] = 32'hFFFFFFF0;
    // rom_array[22308] = 32'hFFFFFFF0;
    // rom_array[22309] = 32'hFFFFFFF1;
    // rom_array[22310] = 32'hFFFFFFF1;
    // rom_array[22311] = 32'hFFFFFFF0;
    // rom_array[22312] = 32'hFFFFFFF0;
    // rom_array[22313] = 32'hFFFFFFF1;
    // rom_array[22314] = 32'hFFFFFFF1;
    // rom_array[22315] = 32'hFFFFFFF0;
    // rom_array[22316] = 32'hFFFFFFF0;
    // rom_array[22317] = 32'hFFFFFFF1;
    // rom_array[22318] = 32'hFFFFFFF1;
    // rom_array[22319] = 32'hFFFFFFF0;
    // rom_array[22320] = 32'hFFFFFFF0;
    // rom_array[22321] = 32'hFFFFFFF1;
    // rom_array[22322] = 32'hFFFFFFF1;
    // rom_array[22323] = 32'hFFFFFFF0;
    // rom_array[22324] = 32'hFFFFFFF0;
    // rom_array[22325] = 32'hFFFFFFF1;
    // rom_array[22326] = 32'hFFFFFFF1;
    // rom_array[22327] = 32'hFFFFFFF0;
    // rom_array[22328] = 32'hFFFFFFF0;
    // rom_array[22329] = 32'hFFFFFFF1;
    // rom_array[22330] = 32'hFFFFFFF1;
    // rom_array[22331] = 32'hFFFFFFF1;
    // rom_array[22332] = 32'hFFFFFFF1;
    // rom_array[22333] = 32'hFFFFFFF1;
    // rom_array[22334] = 32'hFFFFFFF1;
    // rom_array[22335] = 32'hFFFFFFF1;
    // rom_array[22336] = 32'hFFFFFFF1;
    // rom_array[22337] = 32'hFFFFFFF1;
    // rom_array[22338] = 32'hFFFFFFF1;
    // rom_array[22339] = 32'hFFFFFFF1;
    // rom_array[22340] = 32'hFFFFFFF1;
    // rom_array[22341] = 32'hFFFFFFF1;
    // rom_array[22342] = 32'hFFFFFFF1;
    // rom_array[22343] = 32'hFFFFFFF1;
    // rom_array[22344] = 32'hFFFFFFF1;
    // rom_array[22345] = 32'hFFFFFFF1;
    // rom_array[22346] = 32'hFFFFFFF1;
    // rom_array[22347] = 32'hFFFFFFF1;
    // rom_array[22348] = 32'hFFFFFFF1;
    // rom_array[22349] = 32'hFFFFFFF1;
    // rom_array[22350] = 32'hFFFFFFF1;
    // rom_array[22351] = 32'hFFFFFFF1;
    // rom_array[22352] = 32'hFFFFFFF1;
    // rom_array[22353] = 32'hFFFFFFF1;
    // rom_array[22354] = 32'hFFFFFFF1;
    // rom_array[22355] = 32'hFFFFFFF1;
    // rom_array[22356] = 32'hFFFFFFF1;
    // rom_array[22357] = 32'hFFFFFFF1;
    // rom_array[22358] = 32'hFFFFFFF1;
    // rom_array[22359] = 32'hFFFFFFF1;
    // rom_array[22360] = 32'hFFFFFFF1;
    // rom_array[22361] = 32'hFFFFFFF1;
    // rom_array[22362] = 32'hFFFFFFF1;
    // rom_array[22363] = 32'hFFFFFFF1;
    // rom_array[22364] = 32'hFFFFFFF1;
    // rom_array[22365] = 32'hFFFFFFF1;
    // rom_array[22366] = 32'hFFFFFFF1;
    // rom_array[22367] = 32'hFFFFFFF1;
    // rom_array[22368] = 32'hFFFFFFF1;
    // rom_array[22369] = 32'hFFFFFFF1;
    // rom_array[22370] = 32'hFFFFFFF1;
    // rom_array[22371] = 32'hFFFFFFF1;
    // rom_array[22372] = 32'hFFFFFFF1;
    // rom_array[22373] = 32'hFFFFFFF1;
    // rom_array[22374] = 32'hFFFFFFF1;
    // rom_array[22375] = 32'hFFFFFFF1;
    // rom_array[22376] = 32'hFFFFFFF1;
    // rom_array[22377] = 32'hFFFFFFF1;
    // rom_array[22378] = 32'hFFFFFFF1;
    // rom_array[22379] = 32'hFFFFFFF1;
    // rom_array[22380] = 32'hFFFFFFF1;
    // rom_array[22381] = 32'hFFFFFFF1;
    // rom_array[22382] = 32'hFFFFFFF1;
    // rom_array[22383] = 32'hFFFFFFF1;
    // rom_array[22384] = 32'hFFFFFFF1;
    // rom_array[22385] = 32'hFFFFFFF1;
    // rom_array[22386] = 32'hFFFFFFF1;
    // rom_array[22387] = 32'hFFFFFFF1;
    // rom_array[22388] = 32'hFFFFFFF1;
    // rom_array[22389] = 32'hFFFFFFF1;
    // rom_array[22390] = 32'hFFFFFFF1;
    // rom_array[22391] = 32'hFFFFFFF1;
    // rom_array[22392] = 32'hFFFFFFF1;
    // rom_array[22393] = 32'hFFFFFFF1;
    // rom_array[22394] = 32'hFFFFFFF1;
    // rom_array[22395] = 32'hFFFFFFF1;
    // rom_array[22396] = 32'hFFFFFFF1;
    // rom_array[22397] = 32'hFFFFFFF1;
    // rom_array[22398] = 32'hFFFFFFF1;
    // rom_array[22399] = 32'hFFFFFFF1;
    // rom_array[22400] = 32'hFFFFFFF1;
    // rom_array[22401] = 32'hFFFFFFF1;
    // rom_array[22402] = 32'hFFFFFFF1;
    // rom_array[22403] = 32'hFFFFFFF1;
    // rom_array[22404] = 32'hFFFFFFF1;
    // rom_array[22405] = 32'hFFFFFFF1;
    // rom_array[22406] = 32'hFFFFFFF1;
    // rom_array[22407] = 32'hFFFFFFF1;
    // rom_array[22408] = 32'hFFFFFFF1;
    // rom_array[22409] = 32'hFFFFFFF1;
    // rom_array[22410] = 32'hFFFFFFF1;
    // rom_array[22411] = 32'hFFFFFFF1;
    // rom_array[22412] = 32'hFFFFFFF1;
    // rom_array[22413] = 32'hFFFFFFF1;
    // rom_array[22414] = 32'hFFFFFFF1;
    // rom_array[22415] = 32'hFFFFFFF1;
    // rom_array[22416] = 32'hFFFFFFF1;
    // rom_array[22417] = 32'hFFFFFFF1;
    // rom_array[22418] = 32'hFFFFFFF1;
    // rom_array[22419] = 32'hFFFFFFF1;
    // rom_array[22420] = 32'hFFFFFFF1;
    // rom_array[22421] = 32'hFFFFFFF1;
    // rom_array[22422] = 32'hFFFFFFF1;
    // rom_array[22423] = 32'hFFFFFFF1;
    // rom_array[22424] = 32'hFFFFFFF1;
    // rom_array[22425] = 32'hFFFFFFF1;
    // rom_array[22426] = 32'hFFFFFFF1;
    // rom_array[22427] = 32'hFFFFFFF1;
    // rom_array[22428] = 32'hFFFFFFF1;
    // rom_array[22429] = 32'hFFFFFFF1;
    // rom_array[22430] = 32'hFFFFFFF1;
    // rom_array[22431] = 32'hFFFFFFF1;
    // rom_array[22432] = 32'hFFFFFFF1;
    // rom_array[22433] = 32'hFFFFFFF1;
    // rom_array[22434] = 32'hFFFFFFF1;
    // rom_array[22435] = 32'hFFFFFFF1;
    // rom_array[22436] = 32'hFFFFFFF1;
    // rom_array[22437] = 32'hFFFFFFF1;
    // rom_array[22438] = 32'hFFFFFFF1;
    // rom_array[22439] = 32'hFFFFFFF1;
    // rom_array[22440] = 32'hFFFFFFF1;
    // rom_array[22441] = 32'hFFFFFFF1;
    // rom_array[22442] = 32'hFFFFFFF1;
    // rom_array[22443] = 32'hFFFFFFF1;
    // rom_array[22444] = 32'hFFFFFFF1;
    // rom_array[22445] = 32'hFFFFFFF1;
    // rom_array[22446] = 32'hFFFFFFF1;
    // rom_array[22447] = 32'hFFFFFFF1;
    // rom_array[22448] = 32'hFFFFFFF1;
    // rom_array[22449] = 32'hFFFFFFF1;
    // rom_array[22450] = 32'hFFFFFFF1;
    // rom_array[22451] = 32'hFFFFFFF1;
    // rom_array[22452] = 32'hFFFFFFF1;
    // rom_array[22453] = 32'hFFFFFFF1;
    // rom_array[22454] = 32'hFFFFFFF1;
    // rom_array[22455] = 32'hFFFFFFF1;
    // rom_array[22456] = 32'hFFFFFFF1;
    // rom_array[22457] = 32'hFFFFFFF1;
    // rom_array[22458] = 32'hFFFFFFF1;
    // rom_array[22459] = 32'hFFFFFFF1;
    // rom_array[22460] = 32'hFFFFFFF1;
    // rom_array[22461] = 32'hFFFFFFF1;
    // rom_array[22462] = 32'hFFFFFFF1;
    // rom_array[22463] = 32'hFFFFFFF1;
    // rom_array[22464] = 32'hFFFFFFF1;
    // rom_array[22465] = 32'hFFFFFFF1;
    // rom_array[22466] = 32'hFFFFFFF1;
    // rom_array[22467] = 32'hFFFFFFF1;
    // rom_array[22468] = 32'hFFFFFFF1;
    // rom_array[22469] = 32'hFFFFFFF1;
    // rom_array[22470] = 32'hFFFFFFF1;
    // rom_array[22471] = 32'hFFFFFFF1;
    // rom_array[22472] = 32'hFFFFFFF1;
    // rom_array[22473] = 32'hFFFFFFF1;
    // rom_array[22474] = 32'hFFFFFFF1;
    // rom_array[22475] = 32'hFFFFFFF1;
    // rom_array[22476] = 32'hFFFFFFF1;
    // rom_array[22477] = 32'hFFFFFFF1;
    // rom_array[22478] = 32'hFFFFFFF1;
    // rom_array[22479] = 32'hFFFFFFF1;
    // rom_array[22480] = 32'hFFFFFFF1;
    // rom_array[22481] = 32'hFFFFFFF1;
    // rom_array[22482] = 32'hFFFFFFF1;
    // rom_array[22483] = 32'hFFFFFFF1;
    // rom_array[22484] = 32'hFFFFFFF1;
    // rom_array[22485] = 32'hFFFFFFF1;
    // rom_array[22486] = 32'hFFFFFFF1;
    // rom_array[22487] = 32'hFFFFFFF1;
    // rom_array[22488] = 32'hFFFFFFF1;
    // rom_array[22489] = 32'hFFFFFFF1;
    // rom_array[22490] = 32'hFFFFFFF1;
    // rom_array[22491] = 32'hFFFFFFF1;
    // rom_array[22492] = 32'hFFFFFFF1;
    // rom_array[22493] = 32'hFFFFFFF1;
    // rom_array[22494] = 32'hFFFFFFF1;
    // rom_array[22495] = 32'hFFFFFFF1;
    // rom_array[22496] = 32'hFFFFFFF1;
    // rom_array[22497] = 32'hFFFFFFF1;
    // rom_array[22498] = 32'hFFFFFFF1;
    // rom_array[22499] = 32'hFFFFFFF1;
    // rom_array[22500] = 32'hFFFFFFF1;
    // rom_array[22501] = 32'hFFFFFFF1;
    // rom_array[22502] = 32'hFFFFFFF1;
    // rom_array[22503] = 32'hFFFFFFF1;
    // rom_array[22504] = 32'hFFFFFFF1;
    // rom_array[22505] = 32'hFFFFFFF1;
    // rom_array[22506] = 32'hFFFFFFF1;
    // rom_array[22507] = 32'hFFFFFFF1;
    // rom_array[22508] = 32'hFFFFFFF1;
    // rom_array[22509] = 32'hFFFFFFF1;
    // rom_array[22510] = 32'hFFFFFFF1;
    // rom_array[22511] = 32'hFFFFFFF1;
    // rom_array[22512] = 32'hFFFFFFF1;
    // rom_array[22513] = 32'hFFFFFFF1;
    // rom_array[22514] = 32'hFFFFFFF1;
    // rom_array[22515] = 32'hFFFFFFF1;
    // rom_array[22516] = 32'hFFFFFFF1;
    // rom_array[22517] = 32'hFFFFFFF1;
    // rom_array[22518] = 32'hFFFFFFF1;
    // rom_array[22519] = 32'hFFFFFFF1;
    // rom_array[22520] = 32'hFFFFFFF1;
    // rom_array[22521] = 32'hFFFFFFF1;
    // rom_array[22522] = 32'hFFFFFFF1;
    // rom_array[22523] = 32'hFFFFFFF1;
    // rom_array[22524] = 32'hFFFFFFF1;
    // rom_array[22525] = 32'hFFFFFFF1;
    // rom_array[22526] = 32'hFFFFFFF1;
    // rom_array[22527] = 32'hFFFFFFF1;
    // rom_array[22528] = 32'hFFFFFFF1;
    // rom_array[22529] = 32'hFFFFFFF1;
    // rom_array[22530] = 32'hFFFFFFF1;
    // rom_array[22531] = 32'hFFFFFFF1;
    // rom_array[22532] = 32'hFFFFFFF1;
    // rom_array[22533] = 32'hFFFFFFF1;
    // rom_array[22534] = 32'hFFFFFFF1;
    // rom_array[22535] = 32'hFFFFFFF1;
    // rom_array[22536] = 32'hFFFFFFF1;
    // rom_array[22537] = 32'hFFFFFFF1;
    // rom_array[22538] = 32'hFFFFFFF1;
    // rom_array[22539] = 32'hFFFFFFF1;
    // rom_array[22540] = 32'hFFFFFFF1;
    // rom_array[22541] = 32'hFFFFFFF1;
    // rom_array[22542] = 32'hFFFFFFF1;
    // rom_array[22543] = 32'hFFFFFFF1;
    // rom_array[22544] = 32'hFFFFFFF1;
    // rom_array[22545] = 32'hFFFFFFF1;
    // rom_array[22546] = 32'hFFFFFFF1;
    // rom_array[22547] = 32'hFFFFFFF1;
    // rom_array[22548] = 32'hFFFFFFF1;
    // rom_array[22549] = 32'hFFFFFFF1;
    // rom_array[22550] = 32'hFFFFFFF1;
    // rom_array[22551] = 32'hFFFFFFF1;
    // rom_array[22552] = 32'hFFFFFFF1;
    // rom_array[22553] = 32'hFFFFFFF1;
    // rom_array[22554] = 32'hFFFFFFF1;
    // rom_array[22555] = 32'hFFFFFFF1;
    // rom_array[22556] = 32'hFFFFFFF1;
    // rom_array[22557] = 32'hFFFFFFF1;
    // rom_array[22558] = 32'hFFFFFFF1;
    // rom_array[22559] = 32'hFFFFFFF1;
    // rom_array[22560] = 32'hFFFFFFF1;
    // rom_array[22561] = 32'hFFFFFFF1;
    // rom_array[22562] = 32'hFFFFFFF1;
    // rom_array[22563] = 32'hFFFFFFF1;
    // rom_array[22564] = 32'hFFFFFFF1;
    // rom_array[22565] = 32'hFFFFFFF1;
    // rom_array[22566] = 32'hFFFFFFF1;
    // rom_array[22567] = 32'hFFFFFFF1;
    // rom_array[22568] = 32'hFFFFFFF1;
    // rom_array[22569] = 32'hFFFFFFF1;
    // rom_array[22570] = 32'hFFFFFFF1;
    // rom_array[22571] = 32'hFFFFFFF1;
    // rom_array[22572] = 32'hFFFFFFF1;
    // rom_array[22573] = 32'hFFFFFFF1;
    // rom_array[22574] = 32'hFFFFFFF1;
    // rom_array[22575] = 32'hFFFFFFF1;
    // rom_array[22576] = 32'hFFFFFFF1;
    // rom_array[22577] = 32'hFFFFFFF1;
    // rom_array[22578] = 32'hFFFFFFF1;
    // rom_array[22579] = 32'hFFFFFFF1;
    // rom_array[22580] = 32'hFFFFFFF1;
    // rom_array[22581] = 32'hFFFFFFF1;
    // rom_array[22582] = 32'hFFFFFFF1;
    // rom_array[22583] = 32'hFFFFFFF1;
    // rom_array[22584] = 32'hFFFFFFF1;
    // rom_array[22585] = 32'hFFFFFFF1;
    // rom_array[22586] = 32'hFFFFFFF1;
    // rom_array[22587] = 32'hFFFFFFF1;
    // rom_array[22588] = 32'hFFFFFFF1;
    // rom_array[22589] = 32'hFFFFFFF1;
    // rom_array[22590] = 32'hFFFFFFF1;
    // rom_array[22591] = 32'hFFFFFFF1;
    // rom_array[22592] = 32'hFFFFFFF1;
    // rom_array[22593] = 32'hFFFFFFF1;
    // rom_array[22594] = 32'hFFFFFFF1;
    // rom_array[22595] = 32'hFFFFFFF1;
    // rom_array[22596] = 32'hFFFFFFF1;
    // rom_array[22597] = 32'hFFFFFFF1;
    // rom_array[22598] = 32'hFFFFFFF1;
    // rom_array[22599] = 32'hFFFFFFF1;
    // rom_array[22600] = 32'hFFFFFFF1;
    // rom_array[22601] = 32'hFFFFFFF1;
    // rom_array[22602] = 32'hFFFFFFF1;
    // rom_array[22603] = 32'hFFFFFFF1;
    // rom_array[22604] = 32'hFFFFFFF1;
    // rom_array[22605] = 32'hFFFFFFF1;
    // rom_array[22606] = 32'hFFFFFFF1;
    // rom_array[22607] = 32'hFFFFFFF1;
    // rom_array[22608] = 32'hFFFFFFF1;
    // rom_array[22609] = 32'hFFFFFFF1;
    // rom_array[22610] = 32'hFFFFFFF1;
    // rom_array[22611] = 32'hFFFFFFF1;
    // rom_array[22612] = 32'hFFFFFFF1;
    // rom_array[22613] = 32'hFFFFFFF1;
    // rom_array[22614] = 32'hFFFFFFF1;
    // rom_array[22615] = 32'hFFFFFFF1;
    // rom_array[22616] = 32'hFFFFFFF1;
    // rom_array[22617] = 32'hFFFFFFF1;
    // rom_array[22618] = 32'hFFFFFFF1;
    // rom_array[22619] = 32'hFFFFFFF1;
    // rom_array[22620] = 32'hFFFFFFF1;
    // rom_array[22621] = 32'hFFFFFFF1;
    // rom_array[22622] = 32'hFFFFFFF1;
    // rom_array[22623] = 32'hFFFFFFF1;
    // rom_array[22624] = 32'hFFFFFFF1;
    // rom_array[22625] = 32'hFFFFFFF1;
    // rom_array[22626] = 32'hFFFFFFF1;
    // rom_array[22627] = 32'hFFFFFFF1;
    // rom_array[22628] = 32'hFFFFFFF1;
    // rom_array[22629] = 32'hFFFFFFF1;
    // rom_array[22630] = 32'hFFFFFFF1;
    // rom_array[22631] = 32'hFFFFFFF1;
    // rom_array[22632] = 32'hFFFFFFF1;
    // rom_array[22633] = 32'hFFFFFFF1;
    // rom_array[22634] = 32'hFFFFFFF1;
    // rom_array[22635] = 32'hFFFFFFF0;
    // rom_array[22636] = 32'hFFFFFFF0;
    // rom_array[22637] = 32'hFFFFFFF1;
    // rom_array[22638] = 32'hFFFFFFF1;
    // rom_array[22639] = 32'hFFFFFFF0;
    // rom_array[22640] = 32'hFFFFFFF0;
    // rom_array[22641] = 32'hFFFFFFF1;
    // rom_array[22642] = 32'hFFFFFFF1;
    // rom_array[22643] = 32'hFFFFFFF0;
    // rom_array[22644] = 32'hFFFFFFF0;
    // rom_array[22645] = 32'hFFFFFFF1;
    // rom_array[22646] = 32'hFFFFFFF1;
    // rom_array[22647] = 32'hFFFFFFF0;
    // rom_array[22648] = 32'hFFFFFFF0;
    // rom_array[22649] = 32'hFFFFFFF1;
    // rom_array[22650] = 32'hFFFFFFF1;
    // rom_array[22651] = 32'hFFFFFFF0;
    // rom_array[22652] = 32'hFFFFFFF0;
    // rom_array[22653] = 32'hFFFFFFF1;
    // rom_array[22654] = 32'hFFFFFFF1;
    // rom_array[22655] = 32'hFFFFFFF0;
    // rom_array[22656] = 32'hFFFFFFF0;
    // rom_array[22657] = 32'hFFFFFFF1;
    // rom_array[22658] = 32'hFFFFFFF1;
    // rom_array[22659] = 32'hFFFFFFF0;
    // rom_array[22660] = 32'hFFFFFFF0;
    // rom_array[22661] = 32'hFFFFFFF1;
    // rom_array[22662] = 32'hFFFFFFF1;
    // rom_array[22663] = 32'hFFFFFFF0;
    // rom_array[22664] = 32'hFFFFFFF0;
    // rom_array[22665] = 32'hFFFFFFF1;
    // rom_array[22666] = 32'hFFFFFFF1;
    // rom_array[22667] = 32'hFFFFFFF1;
    // rom_array[22668] = 32'hFFFFFFF1;
    // rom_array[22669] = 32'hFFFFFFF1;
    // rom_array[22670] = 32'hFFFFFFF1;
    // rom_array[22671] = 32'hFFFFFFF1;
    // rom_array[22672] = 32'hFFFFFFF1;
    // rom_array[22673] = 32'hFFFFFFF1;
    // rom_array[22674] = 32'hFFFFFFF1;
    // rom_array[22675] = 32'hFFFFFFF1;
    // rom_array[22676] = 32'hFFFFFFF1;
    // rom_array[22677] = 32'hFFFFFFF1;
    // rom_array[22678] = 32'hFFFFFFF1;
    // rom_array[22679] = 32'hFFFFFFF1;
    // rom_array[22680] = 32'hFFFFFFF1;
    // rom_array[22681] = 32'hFFFFFFF1;
    // rom_array[22682] = 32'hFFFFFFF1;
    // rom_array[22683] = 32'hFFFFFFF1;
    // rom_array[22684] = 32'hFFFFFFF1;
    // rom_array[22685] = 32'hFFFFFFF1;
    // rom_array[22686] = 32'hFFFFFFF1;
    // rom_array[22687] = 32'hFFFFFFF1;
    // rom_array[22688] = 32'hFFFFFFF1;
    // rom_array[22689] = 32'hFFFFFFF1;
    // rom_array[22690] = 32'hFFFFFFF1;
    // rom_array[22691] = 32'hFFFFFFF1;
    // rom_array[22692] = 32'hFFFFFFF1;
    // rom_array[22693] = 32'hFFFFFFF1;
    // rom_array[22694] = 32'hFFFFFFF1;
    // rom_array[22695] = 32'hFFFFFFF1;
    // rom_array[22696] = 32'hFFFFFFF1;
    // rom_array[22697] = 32'hFFFFFFF1;
    // rom_array[22698] = 32'hFFFFFFF1;
    // rom_array[22699] = 32'hFFFFFFF1;
    // rom_array[22700] = 32'hFFFFFFF1;
    // rom_array[22701] = 32'hFFFFFFF1;
    // rom_array[22702] = 32'hFFFFFFF1;
    // rom_array[22703] = 32'hFFFFFFF1;
    // rom_array[22704] = 32'hFFFFFFF1;
    // rom_array[22705] = 32'hFFFFFFF1;
    // rom_array[22706] = 32'hFFFFFFF1;
    // rom_array[22707] = 32'hFFFFFFF1;
    // rom_array[22708] = 32'hFFFFFFF1;
    // rom_array[22709] = 32'hFFFFFFF1;
    // rom_array[22710] = 32'hFFFFFFF1;
    // rom_array[22711] = 32'hFFFFFFF1;
    // rom_array[22712] = 32'hFFFFFFF1;
    // rom_array[22713] = 32'hFFFFFFF1;
    // rom_array[22714] = 32'hFFFFFFF1;
    // rom_array[22715] = 32'hFFFFFFF0;
    // rom_array[22716] = 32'hFFFFFFF0;
    // rom_array[22717] = 32'hFFFFFFF1;
    // rom_array[22718] = 32'hFFFFFFF1;
    // rom_array[22719] = 32'hFFFFFFF0;
    // rom_array[22720] = 32'hFFFFFFF0;
    // rom_array[22721] = 32'hFFFFFFF1;
    // rom_array[22722] = 32'hFFFFFFF1;
    // rom_array[22723] = 32'hFFFFFFF0;
    // rom_array[22724] = 32'hFFFFFFF0;
    // rom_array[22725] = 32'hFFFFFFF1;
    // rom_array[22726] = 32'hFFFFFFF1;
    // rom_array[22727] = 32'hFFFFFFF0;
    // rom_array[22728] = 32'hFFFFFFF0;
    // rom_array[22729] = 32'hFFFFFFF1;
    // rom_array[22730] = 32'hFFFFFFF1;
    // rom_array[22731] = 32'hFFFFFFF0;
    // rom_array[22732] = 32'hFFFFFFF0;
    // rom_array[22733] = 32'hFFFFFFF1;
    // rom_array[22734] = 32'hFFFFFFF1;
    // rom_array[22735] = 32'hFFFFFFF0;
    // rom_array[22736] = 32'hFFFFFFF0;
    // rom_array[22737] = 32'hFFFFFFF1;
    // rom_array[22738] = 32'hFFFFFFF1;
    // rom_array[22739] = 32'hFFFFFFF0;
    // rom_array[22740] = 32'hFFFFFFF0;
    // rom_array[22741] = 32'hFFFFFFF1;
    // rom_array[22742] = 32'hFFFFFFF1;
    // rom_array[22743] = 32'hFFFFFFF0;
    // rom_array[22744] = 32'hFFFFFFF0;
    // rom_array[22745] = 32'hFFFFFFF1;
    // rom_array[22746] = 32'hFFFFFFF1;
    // rom_array[22747] = 32'hFFFFFFF0;
    // rom_array[22748] = 32'hFFFFFFF0;
    // rom_array[22749] = 32'hFFFFFFF1;
    // rom_array[22750] = 32'hFFFFFFF1;
    // rom_array[22751] = 32'hFFFFFFF0;
    // rom_array[22752] = 32'hFFFFFFF0;
    // rom_array[22753] = 32'hFFFFFFF1;
    // rom_array[22754] = 32'hFFFFFFF1;
    // rom_array[22755] = 32'hFFFFFFF0;
    // rom_array[22756] = 32'hFFFFFFF0;
    // rom_array[22757] = 32'hFFFFFFF1;
    // rom_array[22758] = 32'hFFFFFFF1;
    // rom_array[22759] = 32'hFFFFFFF0;
    // rom_array[22760] = 32'hFFFFFFF0;
    // rom_array[22761] = 32'hFFFFFFF1;
    // rom_array[22762] = 32'hFFFFFFF1;
    // rom_array[22763] = 32'hFFFFFFF0;
    // rom_array[22764] = 32'hFFFFFFF0;
    // rom_array[22765] = 32'hFFFFFFF1;
    // rom_array[22766] = 32'hFFFFFFF1;
    // rom_array[22767] = 32'hFFFFFFF0;
    // rom_array[22768] = 32'hFFFFFFF0;
    // rom_array[22769] = 32'hFFFFFFF1;
    // rom_array[22770] = 32'hFFFFFFF1;
    // rom_array[22771] = 32'hFFFFFFF0;
    // rom_array[22772] = 32'hFFFFFFF0;
    // rom_array[22773] = 32'hFFFFFFF1;
    // rom_array[22774] = 32'hFFFFFFF1;
    // rom_array[22775] = 32'hFFFFFFF0;
    // rom_array[22776] = 32'hFFFFFFF0;
    // rom_array[22777] = 32'hFFFFFFF1;
    // rom_array[22778] = 32'hFFFFFFF1;
    // rom_array[22779] = 32'hFFFFFFF0;
    // rom_array[22780] = 32'hFFFFFFF0;
    // rom_array[22781] = 32'hFFFFFFF1;
    // rom_array[22782] = 32'hFFFFFFF1;
    // rom_array[22783] = 32'hFFFFFFF0;
    // rom_array[22784] = 32'hFFFFFFF0;
    // rom_array[22785] = 32'hFFFFFFF1;
    // rom_array[22786] = 32'hFFFFFFF1;
    // rom_array[22787] = 32'hFFFFFFF0;
    // rom_array[22788] = 32'hFFFFFFF0;
    // rom_array[22789] = 32'hFFFFFFF1;
    // rom_array[22790] = 32'hFFFFFFF1;
    // rom_array[22791] = 32'hFFFFFFF0;
    // rom_array[22792] = 32'hFFFFFFF0;
    // rom_array[22793] = 32'hFFFFFFF1;
    // rom_array[22794] = 32'hFFFFFFF1;
    // rom_array[22795] = 32'hFFFFFFF0;
    // rom_array[22796] = 32'hFFFFFFF0;
    // rom_array[22797] = 32'hFFFFFFF1;
    // rom_array[22798] = 32'hFFFFFFF1;
    // rom_array[22799] = 32'hFFFFFFF0;
    // rom_array[22800] = 32'hFFFFFFF0;
    // rom_array[22801] = 32'hFFFFFFF1;
    // rom_array[22802] = 32'hFFFFFFF1;
    // rom_array[22803] = 32'hFFFFFFF0;
    // rom_array[22804] = 32'hFFFFFFF0;
    // rom_array[22805] = 32'hFFFFFFF1;
    // rom_array[22806] = 32'hFFFFFFF1;
    // rom_array[22807] = 32'hFFFFFFF0;
    // rom_array[22808] = 32'hFFFFFFF0;
    // rom_array[22809] = 32'hFFFFFFF0;
    // rom_array[22810] = 32'hFFFFFFF0;
    // rom_array[22811] = 32'hFFFFFFF0;
    // rom_array[22812] = 32'hFFFFFFF0;
    // rom_array[22813] = 32'hFFFFFFF1;
    // rom_array[22814] = 32'hFFFFFFF1;
    // rom_array[22815] = 32'hFFFFFFF1;
    // rom_array[22816] = 32'hFFFFFFF1;
    // rom_array[22817] = 32'hFFFFFFF0;
    // rom_array[22818] = 32'hFFFFFFF0;
    // rom_array[22819] = 32'hFFFFFFF0;
    // rom_array[22820] = 32'hFFFFFFF0;
    // rom_array[22821] = 32'hFFFFFFF1;
    // rom_array[22822] = 32'hFFFFFFF1;
    // rom_array[22823] = 32'hFFFFFFF1;
    // rom_array[22824] = 32'hFFFFFFF1;
    // rom_array[22825] = 32'hFFFFFFF0;
    // rom_array[22826] = 32'hFFFFFFF0;
    // rom_array[22827] = 32'hFFFFFFF0;
    // rom_array[22828] = 32'hFFFFFFF0;
    // rom_array[22829] = 32'hFFFFFFF1;
    // rom_array[22830] = 32'hFFFFFFF1;
    // rom_array[22831] = 32'hFFFFFFF1;
    // rom_array[22832] = 32'hFFFFFFF1;
    // rom_array[22833] = 32'hFFFFFFF0;
    // rom_array[22834] = 32'hFFFFFFF0;
    // rom_array[22835] = 32'hFFFFFFF0;
    // rom_array[22836] = 32'hFFFFFFF0;
    // rom_array[22837] = 32'hFFFFFFF1;
    // rom_array[22838] = 32'hFFFFFFF1;
    // rom_array[22839] = 32'hFFFFFFF1;
    // rom_array[22840] = 32'hFFFFFFF1;
    // rom_array[22841] = 32'hFFFFFFF0;
    // rom_array[22842] = 32'hFFFFFFF0;
    // rom_array[22843] = 32'hFFFFFFF0;
    // rom_array[22844] = 32'hFFFFFFF0;
    // rom_array[22845] = 32'hFFFFFFF1;
    // rom_array[22846] = 32'hFFFFFFF1;
    // rom_array[22847] = 32'hFFFFFFF1;
    // rom_array[22848] = 32'hFFFFFFF1;
    // rom_array[22849] = 32'hFFFFFFF0;
    // rom_array[22850] = 32'hFFFFFFF0;
    // rom_array[22851] = 32'hFFFFFFF0;
    // rom_array[22852] = 32'hFFFFFFF0;
    // rom_array[22853] = 32'hFFFFFFF1;
    // rom_array[22854] = 32'hFFFFFFF1;
    // rom_array[22855] = 32'hFFFFFFF1;
    // rom_array[22856] = 32'hFFFFFFF1;
    // rom_array[22857] = 32'hFFFFFFF0;
    // rom_array[22858] = 32'hFFFFFFF0;
    // rom_array[22859] = 32'hFFFFFFF0;
    // rom_array[22860] = 32'hFFFFFFF0;
    // rom_array[22861] = 32'hFFFFFFF1;
    // rom_array[22862] = 32'hFFFFFFF1;
    // rom_array[22863] = 32'hFFFFFFF1;
    // rom_array[22864] = 32'hFFFFFFF1;
    // rom_array[22865] = 32'hFFFFFFF0;
    // rom_array[22866] = 32'hFFFFFFF0;
    // rom_array[22867] = 32'hFFFFFFF0;
    // rom_array[22868] = 32'hFFFFFFF0;
    // rom_array[22869] = 32'hFFFFFFF1;
    // rom_array[22870] = 32'hFFFFFFF1;
    // rom_array[22871] = 32'hFFFFFFF1;
    // rom_array[22872] = 32'hFFFFFFF1;
    // rom_array[22873] = 32'hFFFFFFF1;
    // rom_array[22874] = 32'hFFFFFFF1;
    // rom_array[22875] = 32'hFFFFFFF1;
    // rom_array[22876] = 32'hFFFFFFF1;
    // rom_array[22877] = 32'hFFFFFFF1;
    // rom_array[22878] = 32'hFFFFFFF1;
    // rom_array[22879] = 32'hFFFFFFF1;
    // rom_array[22880] = 32'hFFFFFFF1;
    // rom_array[22881] = 32'hFFFFFFF1;
    // rom_array[22882] = 32'hFFFFFFF1;
    // rom_array[22883] = 32'hFFFFFFF1;
    // rom_array[22884] = 32'hFFFFFFF1;
    // rom_array[22885] = 32'hFFFFFFF1;
    // rom_array[22886] = 32'hFFFFFFF1;
    // rom_array[22887] = 32'hFFFFFFF1;
    // rom_array[22888] = 32'hFFFFFFF1;
    // rom_array[22889] = 32'hFFFFFFF1;
    // rom_array[22890] = 32'hFFFFFFF1;
    // rom_array[22891] = 32'hFFFFFFF1;
    // rom_array[22892] = 32'hFFFFFFF1;
    // rom_array[22893] = 32'hFFFFFFF1;
    // rom_array[22894] = 32'hFFFFFFF1;
    // rom_array[22895] = 32'hFFFFFFF1;
    // rom_array[22896] = 32'hFFFFFFF1;
    // rom_array[22897] = 32'hFFFFFFF1;
    // rom_array[22898] = 32'hFFFFFFF1;
    // rom_array[22899] = 32'hFFFFFFF1;
    // rom_array[22900] = 32'hFFFFFFF1;
    // rom_array[22901] = 32'hFFFFFFF1;
    // rom_array[22902] = 32'hFFFFFFF1;
    // rom_array[22903] = 32'hFFFFFFF1;
    // rom_array[22904] = 32'hFFFFFFF1;
    // rom_array[22905] = 32'hFFFFFFF1;
    // rom_array[22906] = 32'hFFFFFFF1;
    // rom_array[22907] = 32'hFFFFFFF1;
    // rom_array[22908] = 32'hFFFFFFF1;
    // rom_array[22909] = 32'hFFFFFFF1;
    // rom_array[22910] = 32'hFFFFFFF1;
    // rom_array[22911] = 32'hFFFFFFF1;
    // rom_array[22912] = 32'hFFFFFFF1;
    // rom_array[22913] = 32'hFFFFFFF1;
    // rom_array[22914] = 32'hFFFFFFF1;
    // rom_array[22915] = 32'hFFFFFFF1;
    // rom_array[22916] = 32'hFFFFFFF1;
    // rom_array[22917] = 32'hFFFFFFF1;
    // rom_array[22918] = 32'hFFFFFFF1;
    // rom_array[22919] = 32'hFFFFFFF1;
    // rom_array[22920] = 32'hFFFFFFF1;
    // rom_array[22921] = 32'hFFFFFFF1;
    // rom_array[22922] = 32'hFFFFFFF1;
    // rom_array[22923] = 32'hFFFFFFF1;
    // rom_array[22924] = 32'hFFFFFFF1;
    // rom_array[22925] = 32'hFFFFFFF1;
    // rom_array[22926] = 32'hFFFFFFF1;
    // rom_array[22927] = 32'hFFFFFFF1;
    // rom_array[22928] = 32'hFFFFFFF1;
    // rom_array[22929] = 32'hFFFFFFF1;
    // rom_array[22930] = 32'hFFFFFFF1;
    // rom_array[22931] = 32'hFFFFFFF1;
    // rom_array[22932] = 32'hFFFFFFF1;
    // rom_array[22933] = 32'hFFFFFFF1;
    // rom_array[22934] = 32'hFFFFFFF1;
    // rom_array[22935] = 32'hFFFFFFF1;
    // rom_array[22936] = 32'hFFFFFFF1;
    // rom_array[22937] = 32'hFFFFFFF0;
    // rom_array[22938] = 32'hFFFFFFF0;
    // rom_array[22939] = 32'hFFFFFFF0;
    // rom_array[22940] = 32'hFFFFFFF0;
    // rom_array[22941] = 32'hFFFFFFF1;
    // rom_array[22942] = 32'hFFFFFFF1;
    // rom_array[22943] = 32'hFFFFFFF1;
    // rom_array[22944] = 32'hFFFFFFF1;
    // rom_array[22945] = 32'hFFFFFFF0;
    // rom_array[22946] = 32'hFFFFFFF0;
    // rom_array[22947] = 32'hFFFFFFF0;
    // rom_array[22948] = 32'hFFFFFFF0;
    // rom_array[22949] = 32'hFFFFFFF1;
    // rom_array[22950] = 32'hFFFFFFF1;
    // rom_array[22951] = 32'hFFFFFFF1;
    // rom_array[22952] = 32'hFFFFFFF1;
    // rom_array[22953] = 32'hFFFFFFF0;
    // rom_array[22954] = 32'hFFFFFFF0;
    // rom_array[22955] = 32'hFFFFFFF0;
    // rom_array[22956] = 32'hFFFFFFF0;
    // rom_array[22957] = 32'hFFFFFFF1;
    // rom_array[22958] = 32'hFFFFFFF1;
    // rom_array[22959] = 32'hFFFFFFF1;
    // rom_array[22960] = 32'hFFFFFFF1;
    // rom_array[22961] = 32'hFFFFFFF0;
    // rom_array[22962] = 32'hFFFFFFF0;
    // rom_array[22963] = 32'hFFFFFFF0;
    // rom_array[22964] = 32'hFFFFFFF0;
    // rom_array[22965] = 32'hFFFFFFF1;
    // rom_array[22966] = 32'hFFFFFFF1;
    // rom_array[22967] = 32'hFFFFFFF1;
    // rom_array[22968] = 32'hFFFFFFF1;
    // rom_array[22969] = 32'hFFFFFFF0;
    // rom_array[22970] = 32'hFFFFFFF0;
    // rom_array[22971] = 32'hFFFFFFF0;
    // rom_array[22972] = 32'hFFFFFFF0;
    // rom_array[22973] = 32'hFFFFFFF1;
    // rom_array[22974] = 32'hFFFFFFF1;
    // rom_array[22975] = 32'hFFFFFFF1;
    // rom_array[22976] = 32'hFFFFFFF1;
    // rom_array[22977] = 32'hFFFFFFF0;
    // rom_array[22978] = 32'hFFFFFFF0;
    // rom_array[22979] = 32'hFFFFFFF0;
    // rom_array[22980] = 32'hFFFFFFF0;
    // rom_array[22981] = 32'hFFFFFFF1;
    // rom_array[22982] = 32'hFFFFFFF1;
    // rom_array[22983] = 32'hFFFFFFF1;
    // rom_array[22984] = 32'hFFFFFFF1;
    // rom_array[22985] = 32'hFFFFFFF0;
    // rom_array[22986] = 32'hFFFFFFF0;
    // rom_array[22987] = 32'hFFFFFFF0;
    // rom_array[22988] = 32'hFFFFFFF0;
    // rom_array[22989] = 32'hFFFFFFF1;
    // rom_array[22990] = 32'hFFFFFFF1;
    // rom_array[22991] = 32'hFFFFFFF1;
    // rom_array[22992] = 32'hFFFFFFF1;
    // rom_array[22993] = 32'hFFFFFFF0;
    // rom_array[22994] = 32'hFFFFFFF0;
    // rom_array[22995] = 32'hFFFFFFF0;
    // rom_array[22996] = 32'hFFFFFFF0;
    // rom_array[22997] = 32'hFFFFFFF1;
    // rom_array[22998] = 32'hFFFFFFF1;
    // rom_array[22999] = 32'hFFFFFFF1;
    // rom_array[23000] = 32'hFFFFFFF1;
    // rom_array[23001] = 32'hFFFFFFF1;
    // rom_array[23002] = 32'hFFFFFFF1;
    // rom_array[23003] = 32'hFFFFFFF1;
    // rom_array[23004] = 32'hFFFFFFF1;
    // rom_array[23005] = 32'hFFFFFFF1;
    // rom_array[23006] = 32'hFFFFFFF1;
    // rom_array[23007] = 32'hFFFFFFF1;
    // rom_array[23008] = 32'hFFFFFFF1;
    // rom_array[23009] = 32'hFFFFFFF1;
    // rom_array[23010] = 32'hFFFFFFF1;
    // rom_array[23011] = 32'hFFFFFFF1;
    // rom_array[23012] = 32'hFFFFFFF1;
    // rom_array[23013] = 32'hFFFFFFF1;
    // rom_array[23014] = 32'hFFFFFFF1;
    // rom_array[23015] = 32'hFFFFFFF1;
    // rom_array[23016] = 32'hFFFFFFF1;
    // rom_array[23017] = 32'hFFFFFFF1;
    // rom_array[23018] = 32'hFFFFFFF1;
    // rom_array[23019] = 32'hFFFFFFF1;
    // rom_array[23020] = 32'hFFFFFFF1;
    // rom_array[23021] = 32'hFFFFFFF1;
    // rom_array[23022] = 32'hFFFFFFF1;
    // rom_array[23023] = 32'hFFFFFFF1;
    // rom_array[23024] = 32'hFFFFFFF1;
    // rom_array[23025] = 32'hFFFFFFF1;
    // rom_array[23026] = 32'hFFFFFFF1;
    // rom_array[23027] = 32'hFFFFFFF1;
    // rom_array[23028] = 32'hFFFFFFF1;
    // rom_array[23029] = 32'hFFFFFFF1;
    // rom_array[23030] = 32'hFFFFFFF1;
    // rom_array[23031] = 32'hFFFFFFF1;
    // rom_array[23032] = 32'hFFFFFFF1;
    // rom_array[23033] = 32'hFFFFFFF1;
    // rom_array[23034] = 32'hFFFFFFF1;
    // rom_array[23035] = 32'hFFFFFFF1;
    // rom_array[23036] = 32'hFFFFFFF1;
    // rom_array[23037] = 32'hFFFFFFF1;
    // rom_array[23038] = 32'hFFFFFFF1;
    // rom_array[23039] = 32'hFFFFFFF1;
    // rom_array[23040] = 32'hFFFFFFF1;
    // rom_array[23041] = 32'hFFFFFFF1;
    // rom_array[23042] = 32'hFFFFFFF1;
    // rom_array[23043] = 32'hFFFFFFF1;
    // rom_array[23044] = 32'hFFFFFFF1;
    // rom_array[23045] = 32'hFFFFFFF1;
    // rom_array[23046] = 32'hFFFFFFF1;
    // rom_array[23047] = 32'hFFFFFFF1;
    // rom_array[23048] = 32'hFFFFFFF1;
    // rom_array[23049] = 32'hFFFFFFF1;
    // rom_array[23050] = 32'hFFFFFFF1;
    // rom_array[23051] = 32'hFFFFFFF1;
    // rom_array[23052] = 32'hFFFFFFF1;
    // rom_array[23053] = 32'hFFFFFFF1;
    // rom_array[23054] = 32'hFFFFFFF1;
    // rom_array[23055] = 32'hFFFFFFF1;
    // rom_array[23056] = 32'hFFFFFFF1;
    // rom_array[23057] = 32'hFFFFFFF1;
    // rom_array[23058] = 32'hFFFFFFF1;
    // rom_array[23059] = 32'hFFFFFFF1;
    // rom_array[23060] = 32'hFFFFFFF1;
    // rom_array[23061] = 32'hFFFFFFF1;
    // rom_array[23062] = 32'hFFFFFFF1;
    // rom_array[23063] = 32'hFFFFFFF1;
    // rom_array[23064] = 32'hFFFFFFF1;
    // rom_array[23065] = 32'hFFFFFFF1;
    // rom_array[23066] = 32'hFFFFFFF1;
    // rom_array[23067] = 32'hFFFFFFF1;
    // rom_array[23068] = 32'hFFFFFFF1;
    // rom_array[23069] = 32'hFFFFFFF0;
    // rom_array[23070] = 32'hFFFFFFF0;
    // rom_array[23071] = 32'hFFFFFFF0;
    // rom_array[23072] = 32'hFFFFFFF0;
    // rom_array[23073] = 32'hFFFFFFF1;
    // rom_array[23074] = 32'hFFFFFFF1;
    // rom_array[23075] = 32'hFFFFFFF1;
    // rom_array[23076] = 32'hFFFFFFF1;
    // rom_array[23077] = 32'hFFFFFFF0;
    // rom_array[23078] = 32'hFFFFFFF0;
    // rom_array[23079] = 32'hFFFFFFF0;
    // rom_array[23080] = 32'hFFFFFFF0;
    // rom_array[23081] = 32'hFFFFFFF1;
    // rom_array[23082] = 32'hFFFFFFF1;
    // rom_array[23083] = 32'hFFFFFFF1;
    // rom_array[23084] = 32'hFFFFFFF1;
    // rom_array[23085] = 32'hFFFFFFF0;
    // rom_array[23086] = 32'hFFFFFFF0;
    // rom_array[23087] = 32'hFFFFFFF0;
    // rom_array[23088] = 32'hFFFFFFF0;
    // rom_array[23089] = 32'hFFFFFFF1;
    // rom_array[23090] = 32'hFFFFFFF1;
    // rom_array[23091] = 32'hFFFFFFF1;
    // rom_array[23092] = 32'hFFFFFFF1;
    // rom_array[23093] = 32'hFFFFFFF0;
    // rom_array[23094] = 32'hFFFFFFF0;
    // rom_array[23095] = 32'hFFFFFFF0;
    // rom_array[23096] = 32'hFFFFFFF0;
    // rom_array[23097] = 32'hFFFFFFF1;
    // rom_array[23098] = 32'hFFFFFFF1;
    // rom_array[23099] = 32'hFFFFFFF1;
    // rom_array[23100] = 32'hFFFFFFF1;
    // rom_array[23101] = 32'hFFFFFFF0;
    // rom_array[23102] = 32'hFFFFFFF0;
    // rom_array[23103] = 32'hFFFFFFF0;
    // rom_array[23104] = 32'hFFFFFFF0;
    // rom_array[23105] = 32'hFFFFFFF1;
    // rom_array[23106] = 32'hFFFFFFF1;
    // rom_array[23107] = 32'hFFFFFFF1;
    // rom_array[23108] = 32'hFFFFFFF1;
    // rom_array[23109] = 32'hFFFFFFF0;
    // rom_array[23110] = 32'hFFFFFFF0;
    // rom_array[23111] = 32'hFFFFFFF0;
    // rom_array[23112] = 32'hFFFFFFF0;
    // rom_array[23113] = 32'hFFFFFFF1;
    // rom_array[23114] = 32'hFFFFFFF1;
    // rom_array[23115] = 32'hFFFFFFF1;
    // rom_array[23116] = 32'hFFFFFFF1;
    // rom_array[23117] = 32'hFFFFFFF0;
    // rom_array[23118] = 32'hFFFFFFF0;
    // rom_array[23119] = 32'hFFFFFFF0;
    // rom_array[23120] = 32'hFFFFFFF0;
    // rom_array[23121] = 32'hFFFFFFF1;
    // rom_array[23122] = 32'hFFFFFFF1;
    // rom_array[23123] = 32'hFFFFFFF1;
    // rom_array[23124] = 32'hFFFFFFF1;
    // rom_array[23125] = 32'hFFFFFFF0;
    // rom_array[23126] = 32'hFFFFFFF0;
    // rom_array[23127] = 32'hFFFFFFF0;
    // rom_array[23128] = 32'hFFFFFFF0;
    // rom_array[23129] = 32'hFFFFFFF1;
    // rom_array[23130] = 32'hFFFFFFF1;
    // rom_array[23131] = 32'hFFFFFFF1;
    // rom_array[23132] = 32'hFFFFFFF1;
    // rom_array[23133] = 32'hFFFFFFF0;
    // rom_array[23134] = 32'hFFFFFFF0;
    // rom_array[23135] = 32'hFFFFFFF0;
    // rom_array[23136] = 32'hFFFFFFF0;
    // rom_array[23137] = 32'hFFFFFFF1;
    // rom_array[23138] = 32'hFFFFFFF1;
    // rom_array[23139] = 32'hFFFFFFF1;
    // rom_array[23140] = 32'hFFFFFFF1;
    // rom_array[23141] = 32'hFFFFFFF0;
    // rom_array[23142] = 32'hFFFFFFF0;
    // rom_array[23143] = 32'hFFFFFFF0;
    // rom_array[23144] = 32'hFFFFFFF0;
    // rom_array[23145] = 32'hFFFFFFF1;
    // rom_array[23146] = 32'hFFFFFFF1;
    // rom_array[23147] = 32'hFFFFFFF1;
    // rom_array[23148] = 32'hFFFFFFF1;
    // rom_array[23149] = 32'hFFFFFFF0;
    // rom_array[23150] = 32'hFFFFFFF0;
    // rom_array[23151] = 32'hFFFFFFF0;
    // rom_array[23152] = 32'hFFFFFFF0;
    // rom_array[23153] = 32'hFFFFFFF1;
    // rom_array[23154] = 32'hFFFFFFF1;
    // rom_array[23155] = 32'hFFFFFFF1;
    // rom_array[23156] = 32'hFFFFFFF1;
    // rom_array[23157] = 32'hFFFFFFF0;
    // rom_array[23158] = 32'hFFFFFFF0;
    // rom_array[23159] = 32'hFFFFFFF0;
    // rom_array[23160] = 32'hFFFFFFF0;
    // rom_array[23161] = 32'hFFFFFFF1;
    // rom_array[23162] = 32'hFFFFFFF1;
    // rom_array[23163] = 32'hFFFFFFF1;
    // rom_array[23164] = 32'hFFFFFFF1;
    // rom_array[23165] = 32'hFFFFFFF0;
    // rom_array[23166] = 32'hFFFFFFF0;
    // rom_array[23167] = 32'hFFFFFFF0;
    // rom_array[23168] = 32'hFFFFFFF0;
    // rom_array[23169] = 32'hFFFFFFF1;
    // rom_array[23170] = 32'hFFFFFFF1;
    // rom_array[23171] = 32'hFFFFFFF1;
    // rom_array[23172] = 32'hFFFFFFF1;
    // rom_array[23173] = 32'hFFFFFFF0;
    // rom_array[23174] = 32'hFFFFFFF0;
    // rom_array[23175] = 32'hFFFFFFF0;
    // rom_array[23176] = 32'hFFFFFFF0;
    // rom_array[23177] = 32'hFFFFFFF1;
    // rom_array[23178] = 32'hFFFFFFF1;
    // rom_array[23179] = 32'hFFFFFFF1;
    // rom_array[23180] = 32'hFFFFFFF1;
    // rom_array[23181] = 32'hFFFFFFF0;
    // rom_array[23182] = 32'hFFFFFFF0;
    // rom_array[23183] = 32'hFFFFFFF0;
    // rom_array[23184] = 32'hFFFFFFF0;
    // rom_array[23185] = 32'hFFFFFFF1;
    // rom_array[23186] = 32'hFFFFFFF1;
    // rom_array[23187] = 32'hFFFFFFF1;
    // rom_array[23188] = 32'hFFFFFFF1;
    // rom_array[23189] = 32'hFFFFFFF0;
    // rom_array[23190] = 32'hFFFFFFF0;
    // rom_array[23191] = 32'hFFFFFFF0;
    // rom_array[23192] = 32'hFFFFFFF0;
    // rom_array[23193] = 32'hFFFFFFF0;
    // rom_array[23194] = 32'hFFFFFFF0;
    // rom_array[23195] = 32'hFFFFFFF0;
    // rom_array[23196] = 32'hFFFFFFF0;
    // rom_array[23197] = 32'hFFFFFFF1;
    // rom_array[23198] = 32'hFFFFFFF1;
    // rom_array[23199] = 32'hFFFFFFF1;
    // rom_array[23200] = 32'hFFFFFFF1;
    // rom_array[23201] = 32'hFFFFFFF0;
    // rom_array[23202] = 32'hFFFFFFF0;
    // rom_array[23203] = 32'hFFFFFFF0;
    // rom_array[23204] = 32'hFFFFFFF0;
    // rom_array[23205] = 32'hFFFFFFF1;
    // rom_array[23206] = 32'hFFFFFFF1;
    // rom_array[23207] = 32'hFFFFFFF1;
    // rom_array[23208] = 32'hFFFFFFF1;
    // rom_array[23209] = 32'hFFFFFFF0;
    // rom_array[23210] = 32'hFFFFFFF0;
    // rom_array[23211] = 32'hFFFFFFF0;
    // rom_array[23212] = 32'hFFFFFFF0;
    // rom_array[23213] = 32'hFFFFFFF1;
    // rom_array[23214] = 32'hFFFFFFF1;
    // rom_array[23215] = 32'hFFFFFFF1;
    // rom_array[23216] = 32'hFFFFFFF1;
    // rom_array[23217] = 32'hFFFFFFF0;
    // rom_array[23218] = 32'hFFFFFFF0;
    // rom_array[23219] = 32'hFFFFFFF0;
    // rom_array[23220] = 32'hFFFFFFF0;
    // rom_array[23221] = 32'hFFFFFFF1;
    // rom_array[23222] = 32'hFFFFFFF1;
    // rom_array[23223] = 32'hFFFFFFF1;
    // rom_array[23224] = 32'hFFFFFFF1;
    // rom_array[23225] = 32'hFFFFFFF0;
    // rom_array[23226] = 32'hFFFFFFF0;
    // rom_array[23227] = 32'hFFFFFFF0;
    // rom_array[23228] = 32'hFFFFFFF0;
    // rom_array[23229] = 32'hFFFFFFF1;
    // rom_array[23230] = 32'hFFFFFFF1;
    // rom_array[23231] = 32'hFFFFFFF1;
    // rom_array[23232] = 32'hFFFFFFF1;
    // rom_array[23233] = 32'hFFFFFFF0;
    // rom_array[23234] = 32'hFFFFFFF0;
    // rom_array[23235] = 32'hFFFFFFF0;
    // rom_array[23236] = 32'hFFFFFFF0;
    // rom_array[23237] = 32'hFFFFFFF1;
    // rom_array[23238] = 32'hFFFFFFF1;
    // rom_array[23239] = 32'hFFFFFFF1;
    // rom_array[23240] = 32'hFFFFFFF1;
    // rom_array[23241] = 32'hFFFFFFF1;
    // rom_array[23242] = 32'hFFFFFFF1;
    // rom_array[23243] = 32'hFFFFFFF0;
    // rom_array[23244] = 32'hFFFFFFF0;
    // rom_array[23245] = 32'hFFFFFFF1;
    // rom_array[23246] = 32'hFFFFFFF1;
    // rom_array[23247] = 32'hFFFFFFF0;
    // rom_array[23248] = 32'hFFFFFFF0;
    // rom_array[23249] = 32'hFFFFFFF1;
    // rom_array[23250] = 32'hFFFFFFF1;
    // rom_array[23251] = 32'hFFFFFFF0;
    // rom_array[23252] = 32'hFFFFFFF0;
    // rom_array[23253] = 32'hFFFFFFF1;
    // rom_array[23254] = 32'hFFFFFFF1;
    // rom_array[23255] = 32'hFFFFFFF0;
    // rom_array[23256] = 32'hFFFFFFF0;
    // rom_array[23257] = 32'hFFFFFFF1;
    // rom_array[23258] = 32'hFFFFFFF1;
    // rom_array[23259] = 32'hFFFFFFF1;
    // rom_array[23260] = 32'hFFFFFFF1;
    // rom_array[23261] = 32'hFFFFFFF1;
    // rom_array[23262] = 32'hFFFFFFF1;
    // rom_array[23263] = 32'hFFFFFFF1;
    // rom_array[23264] = 32'hFFFFFFF1;
    // rom_array[23265] = 32'hFFFFFFF1;
    // rom_array[23266] = 32'hFFFFFFF1;
    // rom_array[23267] = 32'hFFFFFFF1;
    // rom_array[23268] = 32'hFFFFFFF1;
    // rom_array[23269] = 32'hFFFFFFF1;
    // rom_array[23270] = 32'hFFFFFFF1;
    // rom_array[23271] = 32'hFFFFFFF1;
    // rom_array[23272] = 32'hFFFFFFF1;
    // rom_array[23273] = 32'hFFFFFFF1;
    // rom_array[23274] = 32'hFFFFFFF1;
    // rom_array[23275] = 32'hFFFFFFF0;
    // rom_array[23276] = 32'hFFFFFFF0;
    // rom_array[23277] = 32'hFFFFFFF1;
    // rom_array[23278] = 32'hFFFFFFF1;
    // rom_array[23279] = 32'hFFFFFFF0;
    // rom_array[23280] = 32'hFFFFFFF0;
    // rom_array[23281] = 32'hFFFFFFF1;
    // rom_array[23282] = 32'hFFFFFFF1;
    // rom_array[23283] = 32'hFFFFFFF0;
    // rom_array[23284] = 32'hFFFFFFF0;
    // rom_array[23285] = 32'hFFFFFFF1;
    // rom_array[23286] = 32'hFFFFFFF1;
    // rom_array[23287] = 32'hFFFFFFF0;
    // rom_array[23288] = 32'hFFFFFFF0;
    // rom_array[23289] = 32'hFFFFFFF1;
    // rom_array[23290] = 32'hFFFFFFF1;
    // rom_array[23291] = 32'hFFFFFFF1;
    // rom_array[23292] = 32'hFFFFFFF1;
    // rom_array[23293] = 32'hFFFFFFF1;
    // rom_array[23294] = 32'hFFFFFFF1;
    // rom_array[23295] = 32'hFFFFFFF1;
    // rom_array[23296] = 32'hFFFFFFF1;
    // rom_array[23297] = 32'hFFFFFFF1;
    // rom_array[23298] = 32'hFFFFFFF1;
    // rom_array[23299] = 32'hFFFFFFF1;
    // rom_array[23300] = 32'hFFFFFFF1;
    // rom_array[23301] = 32'hFFFFFFF1;
    // rom_array[23302] = 32'hFFFFFFF1;
    // rom_array[23303] = 32'hFFFFFFF1;
    // rom_array[23304] = 32'hFFFFFFF1;
    // rom_array[23305] = 32'hFFFFFFF1;
    // rom_array[23306] = 32'hFFFFFFF1;
    // rom_array[23307] = 32'hFFFFFFF1;
    // rom_array[23308] = 32'hFFFFFFF1;
    // rom_array[23309] = 32'hFFFFFFF1;
    // rom_array[23310] = 32'hFFFFFFF1;
    // rom_array[23311] = 32'hFFFFFFF1;
    // rom_array[23312] = 32'hFFFFFFF1;
    // rom_array[23313] = 32'hFFFFFFF1;
    // rom_array[23314] = 32'hFFFFFFF1;
    // rom_array[23315] = 32'hFFFFFFF1;
    // rom_array[23316] = 32'hFFFFFFF1;
    // rom_array[23317] = 32'hFFFFFFF1;
    // rom_array[23318] = 32'hFFFFFFF1;
    // rom_array[23319] = 32'hFFFFFFF1;
    // rom_array[23320] = 32'hFFFFFFF1;
    // rom_array[23321] = 32'hFFFFFFF1;
    // rom_array[23322] = 32'hFFFFFFF1;
    // rom_array[23323] = 32'hFFFFFFF1;
    // rom_array[23324] = 32'hFFFFFFF1;
    // rom_array[23325] = 32'hFFFFFFF1;
    // rom_array[23326] = 32'hFFFFFFF1;
    // rom_array[23327] = 32'hFFFFFFF1;
    // rom_array[23328] = 32'hFFFFFFF1;
    // rom_array[23329] = 32'hFFFFFFF1;
    // rom_array[23330] = 32'hFFFFFFF1;
    // rom_array[23331] = 32'hFFFFFFF1;
    // rom_array[23332] = 32'hFFFFFFF1;
    // rom_array[23333] = 32'hFFFFFFF1;
    // rom_array[23334] = 32'hFFFFFFF1;
    // rom_array[23335] = 32'hFFFFFFF1;
    // rom_array[23336] = 32'hFFFFFFF1;
    // rom_array[23337] = 32'hFFFFFFF1;
    // rom_array[23338] = 32'hFFFFFFF1;
    // rom_array[23339] = 32'hFFFFFFF0;
    // rom_array[23340] = 32'hFFFFFFF0;
    // rom_array[23341] = 32'hFFFFFFF1;
    // rom_array[23342] = 32'hFFFFFFF1;
    // rom_array[23343] = 32'hFFFFFFF0;
    // rom_array[23344] = 32'hFFFFFFF0;
    // rom_array[23345] = 32'hFFFFFFF1;
    // rom_array[23346] = 32'hFFFFFFF1;
    // rom_array[23347] = 32'hFFFFFFF0;
    // rom_array[23348] = 32'hFFFFFFF0;
    // rom_array[23349] = 32'hFFFFFFF1;
    // rom_array[23350] = 32'hFFFFFFF1;
    // rom_array[23351] = 32'hFFFFFFF0;
    // rom_array[23352] = 32'hFFFFFFF0;
    // rom_array[23353] = 32'hFFFFFFF1;
    // rom_array[23354] = 32'hFFFFFFF1;
    // rom_array[23355] = 32'hFFFFFFF1;
    // rom_array[23356] = 32'hFFFFFFF1;
    // rom_array[23357] = 32'hFFFFFFF1;
    // rom_array[23358] = 32'hFFFFFFF1;
    // rom_array[23359] = 32'hFFFFFFF1;
    // rom_array[23360] = 32'hFFFFFFF1;
    // rom_array[23361] = 32'hFFFFFFF1;
    // rom_array[23362] = 32'hFFFFFFF1;
    // rom_array[23363] = 32'hFFFFFFF1;
    // rom_array[23364] = 32'hFFFFFFF1;
    // rom_array[23365] = 32'hFFFFFFF1;
    // rom_array[23366] = 32'hFFFFFFF1;
    // rom_array[23367] = 32'hFFFFFFF1;
    // rom_array[23368] = 32'hFFFFFFF1;
    // rom_array[23369] = 32'hFFFFFFF1;
    // rom_array[23370] = 32'hFFFFFFF1;
    // rom_array[23371] = 32'hFFFFFFF0;
    // rom_array[23372] = 32'hFFFFFFF0;
    // rom_array[23373] = 32'hFFFFFFF1;
    // rom_array[23374] = 32'hFFFFFFF1;
    // rom_array[23375] = 32'hFFFFFFF0;
    // rom_array[23376] = 32'hFFFFFFF0;
    // rom_array[23377] = 32'hFFFFFFF1;
    // rom_array[23378] = 32'hFFFFFFF1;
    // rom_array[23379] = 32'hFFFFFFF0;
    // rom_array[23380] = 32'hFFFFFFF0;
    // rom_array[23381] = 32'hFFFFFFF1;
    // rom_array[23382] = 32'hFFFFFFF1;
    // rom_array[23383] = 32'hFFFFFFF0;
    // rom_array[23384] = 32'hFFFFFFF0;
    // rom_array[23385] = 32'hFFFFFFF1;
    // rom_array[23386] = 32'hFFFFFFF1;
    // rom_array[23387] = 32'hFFFFFFF1;
    // rom_array[23388] = 32'hFFFFFFF1;
    // rom_array[23389] = 32'hFFFFFFF0;
    // rom_array[23390] = 32'hFFFFFFF0;
    // rom_array[23391] = 32'hFFFFFFF0;
    // rom_array[23392] = 32'hFFFFFFF0;
    // rom_array[23393] = 32'hFFFFFFF1;
    // rom_array[23394] = 32'hFFFFFFF1;
    // rom_array[23395] = 32'hFFFFFFF1;
    // rom_array[23396] = 32'hFFFFFFF1;
    // rom_array[23397] = 32'hFFFFFFF0;
    // rom_array[23398] = 32'hFFFFFFF0;
    // rom_array[23399] = 32'hFFFFFFF0;
    // rom_array[23400] = 32'hFFFFFFF0;
    // rom_array[23401] = 32'hFFFFFFF1;
    // rom_array[23402] = 32'hFFFFFFF1;
    // rom_array[23403] = 32'hFFFFFFF1;
    // rom_array[23404] = 32'hFFFFFFF1;
    // rom_array[23405] = 32'hFFFFFFF0;
    // rom_array[23406] = 32'hFFFFFFF0;
    // rom_array[23407] = 32'hFFFFFFF0;
    // rom_array[23408] = 32'hFFFFFFF0;
    // rom_array[23409] = 32'hFFFFFFF1;
    // rom_array[23410] = 32'hFFFFFFF1;
    // rom_array[23411] = 32'hFFFFFFF1;
    // rom_array[23412] = 32'hFFFFFFF1;
    // rom_array[23413] = 32'hFFFFFFF0;
    // rom_array[23414] = 32'hFFFFFFF0;
    // rom_array[23415] = 32'hFFFFFFF0;
    // rom_array[23416] = 32'hFFFFFFF0;
    // rom_array[23417] = 32'hFFFFFFF1;
    // rom_array[23418] = 32'hFFFFFFF1;
    // rom_array[23419] = 32'hFFFFFFF1;
    // rom_array[23420] = 32'hFFFFFFF1;
    // rom_array[23421] = 32'hFFFFFFF0;
    // rom_array[23422] = 32'hFFFFFFF0;
    // rom_array[23423] = 32'hFFFFFFF0;
    // rom_array[23424] = 32'hFFFFFFF0;
    // rom_array[23425] = 32'hFFFFFFF1;
    // rom_array[23426] = 32'hFFFFFFF1;
    // rom_array[23427] = 32'hFFFFFFF1;
    // rom_array[23428] = 32'hFFFFFFF1;
    // rom_array[23429] = 32'hFFFFFFF0;
    // rom_array[23430] = 32'hFFFFFFF0;
    // rom_array[23431] = 32'hFFFFFFF0;
    // rom_array[23432] = 32'hFFFFFFF0;
    // rom_array[23433] = 32'hFFFFFFF0;
    // rom_array[23434] = 32'hFFFFFFF0;
    // rom_array[23435] = 32'hFFFFFFF0;
    // rom_array[23436] = 32'hFFFFFFF0;
    // rom_array[23437] = 32'hFFFFFFF1;
    // rom_array[23438] = 32'hFFFFFFF1;
    // rom_array[23439] = 32'hFFFFFFF1;
    // rom_array[23440] = 32'hFFFFFFF1;
    // rom_array[23441] = 32'hFFFFFFF0;
    // rom_array[23442] = 32'hFFFFFFF0;
    // rom_array[23443] = 32'hFFFFFFF0;
    // rom_array[23444] = 32'hFFFFFFF0;
    // rom_array[23445] = 32'hFFFFFFF1;
    // rom_array[23446] = 32'hFFFFFFF1;
    // rom_array[23447] = 32'hFFFFFFF1;
    // rom_array[23448] = 32'hFFFFFFF1;
    // rom_array[23449] = 32'hFFFFFFF0;
    // rom_array[23450] = 32'hFFFFFFF0;
    // rom_array[23451] = 32'hFFFFFFF0;
    // rom_array[23452] = 32'hFFFFFFF0;
    // rom_array[23453] = 32'hFFFFFFF1;
    // rom_array[23454] = 32'hFFFFFFF1;
    // rom_array[23455] = 32'hFFFFFFF1;
    // rom_array[23456] = 32'hFFFFFFF1;
    // rom_array[23457] = 32'hFFFFFFF0;
    // rom_array[23458] = 32'hFFFFFFF0;
    // rom_array[23459] = 32'hFFFFFFF0;
    // rom_array[23460] = 32'hFFFFFFF0;
    // rom_array[23461] = 32'hFFFFFFF1;
    // rom_array[23462] = 32'hFFFFFFF1;
    // rom_array[23463] = 32'hFFFFFFF1;
    // rom_array[23464] = 32'hFFFFFFF1;
    // rom_array[23465] = 32'hFFFFFFF0;
    // rom_array[23466] = 32'hFFFFFFF0;
    // rom_array[23467] = 32'hFFFFFFF0;
    // rom_array[23468] = 32'hFFFFFFF0;
    // rom_array[23469] = 32'hFFFFFFF1;
    // rom_array[23470] = 32'hFFFFFFF1;
    // rom_array[23471] = 32'hFFFFFFF1;
    // rom_array[23472] = 32'hFFFFFFF1;
    // rom_array[23473] = 32'hFFFFFFF0;
    // rom_array[23474] = 32'hFFFFFFF0;
    // rom_array[23475] = 32'hFFFFFFF0;
    // rom_array[23476] = 32'hFFFFFFF0;
    // rom_array[23477] = 32'hFFFFFFF1;
    // rom_array[23478] = 32'hFFFFFFF1;
    // rom_array[23479] = 32'hFFFFFFF1;
    // rom_array[23480] = 32'hFFFFFFF1;
    // rom_array[23481] = 32'hFFFFFFF0;
    // rom_array[23482] = 32'hFFFFFFF0;
    // rom_array[23483] = 32'hFFFFFFF0;
    // rom_array[23484] = 32'hFFFFFFF0;
    // rom_array[23485] = 32'hFFFFFFF1;
    // rom_array[23486] = 32'hFFFFFFF1;
    // rom_array[23487] = 32'hFFFFFFF1;
    // rom_array[23488] = 32'hFFFFFFF1;
    // rom_array[23489] = 32'hFFFFFFF0;
    // rom_array[23490] = 32'hFFFFFFF0;
    // rom_array[23491] = 32'hFFFFFFF0;
    // rom_array[23492] = 32'hFFFFFFF0;
    // rom_array[23493] = 32'hFFFFFFF1;
    // rom_array[23494] = 32'hFFFFFFF1;
    // rom_array[23495] = 32'hFFFFFFF1;
    // rom_array[23496] = 32'hFFFFFFF1;
    // rom_array[23497] = 32'hFFFFFFF0;
    // rom_array[23498] = 32'hFFFFFFF0;
    // rom_array[23499] = 32'hFFFFFFF0;
    // rom_array[23500] = 32'hFFFFFFF0;
    // rom_array[23501] = 32'hFFFFFFF1;
    // rom_array[23502] = 32'hFFFFFFF1;
    // rom_array[23503] = 32'hFFFFFFF1;
    // rom_array[23504] = 32'hFFFFFFF1;
    // rom_array[23505] = 32'hFFFFFFF0;
    // rom_array[23506] = 32'hFFFFFFF0;
    // rom_array[23507] = 32'hFFFFFFF0;
    // rom_array[23508] = 32'hFFFFFFF0;
    // rom_array[23509] = 32'hFFFFFFF1;
    // rom_array[23510] = 32'hFFFFFFF1;
    // rom_array[23511] = 32'hFFFFFFF1;
    // rom_array[23512] = 32'hFFFFFFF1;
    // rom_array[23513] = 32'hFFFFFFF0;
    // rom_array[23514] = 32'hFFFFFFF0;
    // rom_array[23515] = 32'hFFFFFFF0;
    // rom_array[23516] = 32'hFFFFFFF0;
    // rom_array[23517] = 32'hFFFFFFF1;
    // rom_array[23518] = 32'hFFFFFFF1;
    // rom_array[23519] = 32'hFFFFFFF1;
    // rom_array[23520] = 32'hFFFFFFF1;
    // rom_array[23521] = 32'hFFFFFFF0;
    // rom_array[23522] = 32'hFFFFFFF0;
    // rom_array[23523] = 32'hFFFFFFF0;
    // rom_array[23524] = 32'hFFFFFFF0;
    // rom_array[23525] = 32'hFFFFFFF1;
    // rom_array[23526] = 32'hFFFFFFF1;
    // rom_array[23527] = 32'hFFFFFFF1;
    // rom_array[23528] = 32'hFFFFFFF1;
    // rom_array[23529] = 32'hFFFFFFF0;
    // rom_array[23530] = 32'hFFFFFFF0;
    // rom_array[23531] = 32'hFFFFFFF0;
    // rom_array[23532] = 32'hFFFFFFF0;
    // rom_array[23533] = 32'hFFFFFFF1;
    // rom_array[23534] = 32'hFFFFFFF1;
    // rom_array[23535] = 32'hFFFFFFF1;
    // rom_array[23536] = 32'hFFFFFFF1;
    // rom_array[23537] = 32'hFFFFFFF0;
    // rom_array[23538] = 32'hFFFFFFF0;
    // rom_array[23539] = 32'hFFFFFFF0;
    // rom_array[23540] = 32'hFFFFFFF0;
    // rom_array[23541] = 32'hFFFFFFF1;
    // rom_array[23542] = 32'hFFFFFFF1;
    // rom_array[23543] = 32'hFFFFFFF1;
    // rom_array[23544] = 32'hFFFFFFF1;
    // rom_array[23545] = 32'hFFFFFFF0;
    // rom_array[23546] = 32'hFFFFFFF0;
    // rom_array[23547] = 32'hFFFFFFF0;
    // rom_array[23548] = 32'hFFFFFFF0;
    // rom_array[23549] = 32'hFFFFFFF1;
    // rom_array[23550] = 32'hFFFFFFF1;
    // rom_array[23551] = 32'hFFFFFFF1;
    // rom_array[23552] = 32'hFFFFFFF1;
    // rom_array[23553] = 32'hFFFFFFF0;
    // rom_array[23554] = 32'hFFFFFFF0;
    // rom_array[23555] = 32'hFFFFFFF0;
    // rom_array[23556] = 32'hFFFFFFF0;
    // rom_array[23557] = 32'hFFFFFFF1;
    // rom_array[23558] = 32'hFFFFFFF1;
    // rom_array[23559] = 32'hFFFFFFF1;
    // rom_array[23560] = 32'hFFFFFFF1;
    // rom_array[23561] = 32'hFFFFFFF1;
    // rom_array[23562] = 32'hFFFFFFF1;
    // rom_array[23563] = 32'hFFFFFFF1;
    // rom_array[23564] = 32'hFFFFFFF1;
    // rom_array[23565] = 32'hFFFFFFF1;
    // rom_array[23566] = 32'hFFFFFFF1;
    // rom_array[23567] = 32'hFFFFFFF1;
    // rom_array[23568] = 32'hFFFFFFF1;
    // rom_array[23569] = 32'hFFFFFFF1;
    // rom_array[23570] = 32'hFFFFFFF1;
    // rom_array[23571] = 32'hFFFFFFF1;
    // rom_array[23572] = 32'hFFFFFFF1;
    // rom_array[23573] = 32'hFFFFFFF1;
    // rom_array[23574] = 32'hFFFFFFF1;
    // rom_array[23575] = 32'hFFFFFFF1;
    // rom_array[23576] = 32'hFFFFFFF1;
    // rom_array[23577] = 32'hFFFFFFF1;
    // rom_array[23578] = 32'hFFFFFFF1;
    // rom_array[23579] = 32'hFFFFFFF1;
    // rom_array[23580] = 32'hFFFFFFF1;
    // rom_array[23581] = 32'hFFFFFFF0;
    // rom_array[23582] = 32'hFFFFFFF0;
    // rom_array[23583] = 32'hFFFFFFF0;
    // rom_array[23584] = 32'hFFFFFFF0;
    // rom_array[23585] = 32'hFFFFFFF1;
    // rom_array[23586] = 32'hFFFFFFF1;
    // rom_array[23587] = 32'hFFFFFFF1;
    // rom_array[23588] = 32'hFFFFFFF1;
    // rom_array[23589] = 32'hFFFFFFF0;
    // rom_array[23590] = 32'hFFFFFFF0;
    // rom_array[23591] = 32'hFFFFFFF0;
    // rom_array[23592] = 32'hFFFFFFF0;
    // rom_array[23593] = 32'hFFFFFFF1;
    // rom_array[23594] = 32'hFFFFFFF1;
    // rom_array[23595] = 32'hFFFFFFF1;
    // rom_array[23596] = 32'hFFFFFFF1;
    // rom_array[23597] = 32'hFFFFFFF1;
    // rom_array[23598] = 32'hFFFFFFF1;
    // rom_array[23599] = 32'hFFFFFFF1;
    // rom_array[23600] = 32'hFFFFFFF1;
    // rom_array[23601] = 32'hFFFFFFF1;
    // rom_array[23602] = 32'hFFFFFFF1;
    // rom_array[23603] = 32'hFFFFFFF1;
    // rom_array[23604] = 32'hFFFFFFF1;
    // rom_array[23605] = 32'hFFFFFFF1;
    // rom_array[23606] = 32'hFFFFFFF1;
    // rom_array[23607] = 32'hFFFFFFF1;
    // rom_array[23608] = 32'hFFFFFFF1;
    // rom_array[23609] = 32'hFFFFFFF1;
    // rom_array[23610] = 32'hFFFFFFF1;
    // rom_array[23611] = 32'hFFFFFFF1;
    // rom_array[23612] = 32'hFFFFFFF1;
    // rom_array[23613] = 32'hFFFFFFF0;
    // rom_array[23614] = 32'hFFFFFFF0;
    // rom_array[23615] = 32'hFFFFFFF0;
    // rom_array[23616] = 32'hFFFFFFF0;
    // rom_array[23617] = 32'hFFFFFFF1;
    // rom_array[23618] = 32'hFFFFFFF1;
    // rom_array[23619] = 32'hFFFFFFF1;
    // rom_array[23620] = 32'hFFFFFFF1;
    // rom_array[23621] = 32'hFFFFFFF0;
    // rom_array[23622] = 32'hFFFFFFF0;
    // rom_array[23623] = 32'hFFFFFFF0;
    // rom_array[23624] = 32'hFFFFFFF0;
    // rom_array[23625] = 32'hFFFFFFF1;
    // rom_array[23626] = 32'hFFFFFFF1;
    // rom_array[23627] = 32'hFFFFFFF1;
    // rom_array[23628] = 32'hFFFFFFF1;
    // rom_array[23629] = 32'hFFFFFFF0;
    // rom_array[23630] = 32'hFFFFFFF0;
    // rom_array[23631] = 32'hFFFFFFF0;
    // rom_array[23632] = 32'hFFFFFFF0;
    // rom_array[23633] = 32'hFFFFFFF1;
    // rom_array[23634] = 32'hFFFFFFF1;
    // rom_array[23635] = 32'hFFFFFFF1;
    // rom_array[23636] = 32'hFFFFFFF1;
    // rom_array[23637] = 32'hFFFFFFF0;
    // rom_array[23638] = 32'hFFFFFFF0;
    // rom_array[23639] = 32'hFFFFFFF0;
    // rom_array[23640] = 32'hFFFFFFF0;
    // rom_array[23641] = 32'hFFFFFFF1;
    // rom_array[23642] = 32'hFFFFFFF1;
    // rom_array[23643] = 32'hFFFFFFF1;
    // rom_array[23644] = 32'hFFFFFFF1;
    // rom_array[23645] = 32'hFFFFFFF1;
    // rom_array[23646] = 32'hFFFFFFF1;
    // rom_array[23647] = 32'hFFFFFFF1;
    // rom_array[23648] = 32'hFFFFFFF1;
    // rom_array[23649] = 32'hFFFFFFF1;
    // rom_array[23650] = 32'hFFFFFFF1;
    // rom_array[23651] = 32'hFFFFFFF1;
    // rom_array[23652] = 32'hFFFFFFF1;
    // rom_array[23653] = 32'hFFFFFFF1;
    // rom_array[23654] = 32'hFFFFFFF1;
    // rom_array[23655] = 32'hFFFFFFF1;
    // rom_array[23656] = 32'hFFFFFFF1;
    // rom_array[23657] = 32'hFFFFFFF1;
    // rom_array[23658] = 32'hFFFFFFF1;
    // rom_array[23659] = 32'hFFFFFFF1;
    // rom_array[23660] = 32'hFFFFFFF1;
    // rom_array[23661] = 32'hFFFFFFF1;
    // rom_array[23662] = 32'hFFFFFFF1;
    // rom_array[23663] = 32'hFFFFFFF1;
    // rom_array[23664] = 32'hFFFFFFF1;
    // rom_array[23665] = 32'hFFFFFFF1;
    // rom_array[23666] = 32'hFFFFFFF1;
    // rom_array[23667] = 32'hFFFFFFF1;
    // rom_array[23668] = 32'hFFFFFFF1;
    // rom_array[23669] = 32'hFFFFFFF1;
    // rom_array[23670] = 32'hFFFFFFF1;
    // rom_array[23671] = 32'hFFFFFFF1;
    // rom_array[23672] = 32'hFFFFFFF1;
    // rom_array[23673] = 32'hFFFFFFF1;
    // rom_array[23674] = 32'hFFFFFFF1;
    // rom_array[23675] = 32'hFFFFFFF1;
    // rom_array[23676] = 32'hFFFFFFF1;
    // rom_array[23677] = 32'hFFFFFFF0;
    // rom_array[23678] = 32'hFFFFFFF0;
    // rom_array[23679] = 32'hFFFFFFF0;
    // rom_array[23680] = 32'hFFFFFFF0;
    // rom_array[23681] = 32'hFFFFFFF1;
    // rom_array[23682] = 32'hFFFFFFF1;
    // rom_array[23683] = 32'hFFFFFFF1;
    // rom_array[23684] = 32'hFFFFFFF1;
    // rom_array[23685] = 32'hFFFFFFF0;
    // rom_array[23686] = 32'hFFFFFFF0;
    // rom_array[23687] = 32'hFFFFFFF0;
    // rom_array[23688] = 32'hFFFFFFF0;
    // rom_array[23689] = 32'hFFFFFFF1;
    // rom_array[23690] = 32'hFFFFFFF1;
    // rom_array[23691] = 32'hFFFFFFF1;
    // rom_array[23692] = 32'hFFFFFFF1;
    // rom_array[23693] = 32'hFFFFFFF0;
    // rom_array[23694] = 32'hFFFFFFF0;
    // rom_array[23695] = 32'hFFFFFFF0;
    // rom_array[23696] = 32'hFFFFFFF0;
    // rom_array[23697] = 32'hFFFFFFF1;
    // rom_array[23698] = 32'hFFFFFFF1;
    // rom_array[23699] = 32'hFFFFFFF1;
    // rom_array[23700] = 32'hFFFFFFF1;
    // rom_array[23701] = 32'hFFFFFFF0;
    // rom_array[23702] = 32'hFFFFFFF0;
    // rom_array[23703] = 32'hFFFFFFF0;
    // rom_array[23704] = 32'hFFFFFFF0;
    // rom_array[23705] = 32'hFFFFFFF1;
    // rom_array[23706] = 32'hFFFFFFF1;
    // rom_array[23707] = 32'hFFFFFFF1;
    // rom_array[23708] = 32'hFFFFFFF1;
    // rom_array[23709] = 32'hFFFFFFF0;
    // rom_array[23710] = 32'hFFFFFFF0;
    // rom_array[23711] = 32'hFFFFFFF1;
    // rom_array[23712] = 32'hFFFFFFF1;
    // rom_array[23713] = 32'hFFFFFFF1;
    // rom_array[23714] = 32'hFFFFFFF1;
    // rom_array[23715] = 32'hFFFFFFF1;
    // rom_array[23716] = 32'hFFFFFFF1;
    // rom_array[23717] = 32'hFFFFFFF0;
    // rom_array[23718] = 32'hFFFFFFF0;
    // rom_array[23719] = 32'hFFFFFFF1;
    // rom_array[23720] = 32'hFFFFFFF1;
    // rom_array[23721] = 32'hFFFFFFF1;
    // rom_array[23722] = 32'hFFFFFFF1;
    // rom_array[23723] = 32'hFFFFFFF1;
    // rom_array[23724] = 32'hFFFFFFF1;
    // rom_array[23725] = 32'hFFFFFFF1;
    // rom_array[23726] = 32'hFFFFFFF1;
    // rom_array[23727] = 32'hFFFFFFF1;
    // rom_array[23728] = 32'hFFFFFFF1;
    // rom_array[23729] = 32'hFFFFFFF1;
    // rom_array[23730] = 32'hFFFFFFF1;
    // rom_array[23731] = 32'hFFFFFFF1;
    // rom_array[23732] = 32'hFFFFFFF1;
    // rom_array[23733] = 32'hFFFFFFF1;
    // rom_array[23734] = 32'hFFFFFFF1;
    // rom_array[23735] = 32'hFFFFFFF1;
    // rom_array[23736] = 32'hFFFFFFF1;
    // rom_array[23737] = 32'hFFFFFFF0;
    // rom_array[23738] = 32'hFFFFFFF0;
    // rom_array[23739] = 32'hFFFFFFF1;
    // rom_array[23740] = 32'hFFFFFFF1;
    // rom_array[23741] = 32'hFFFFFFF0;
    // rom_array[23742] = 32'hFFFFFFF0;
    // rom_array[23743] = 32'hFFFFFFF1;
    // rom_array[23744] = 32'hFFFFFFF1;
    // rom_array[23745] = 32'hFFFFFFF0;
    // rom_array[23746] = 32'hFFFFFFF0;
    // rom_array[23747] = 32'hFFFFFFF1;
    // rom_array[23748] = 32'hFFFFFFF1;
    // rom_array[23749] = 32'hFFFFFFF0;
    // rom_array[23750] = 32'hFFFFFFF0;
    // rom_array[23751] = 32'hFFFFFFF1;
    // rom_array[23752] = 32'hFFFFFFF1;
    // rom_array[23753] = 32'hFFFFFFF0;
    // rom_array[23754] = 32'hFFFFFFF0;
    // rom_array[23755] = 32'hFFFFFFF1;
    // rom_array[23756] = 32'hFFFFFFF1;
    // rom_array[23757] = 32'hFFFFFFF0;
    // rom_array[23758] = 32'hFFFFFFF0;
    // rom_array[23759] = 32'hFFFFFFF1;
    // rom_array[23760] = 32'hFFFFFFF1;
    // rom_array[23761] = 32'hFFFFFFF0;
    // rom_array[23762] = 32'hFFFFFFF0;
    // rom_array[23763] = 32'hFFFFFFF1;
    // rom_array[23764] = 32'hFFFFFFF1;
    // rom_array[23765] = 32'hFFFFFFF0;
    // rom_array[23766] = 32'hFFFFFFF0;
    // rom_array[23767] = 32'hFFFFFFF1;
    // rom_array[23768] = 32'hFFFFFFF1;
    // rom_array[23769] = 32'hFFFFFFF0;
    // rom_array[23770] = 32'hFFFFFFF0;
    // rom_array[23771] = 32'hFFFFFFF1;
    // rom_array[23772] = 32'hFFFFFFF1;
    // rom_array[23773] = 32'hFFFFFFF0;
    // rom_array[23774] = 32'hFFFFFFF0;
    // rom_array[23775] = 32'hFFFFFFF1;
    // rom_array[23776] = 32'hFFFFFFF1;
    // rom_array[23777] = 32'hFFFFFFF0;
    // rom_array[23778] = 32'hFFFFFFF0;
    // rom_array[23779] = 32'hFFFFFFF1;
    // rom_array[23780] = 32'hFFFFFFF1;
    // rom_array[23781] = 32'hFFFFFFF0;
    // rom_array[23782] = 32'hFFFFFFF0;
    // rom_array[23783] = 32'hFFFFFFF1;
    // rom_array[23784] = 32'hFFFFFFF1;
    // rom_array[23785] = 32'hFFFFFFF0;
    // rom_array[23786] = 32'hFFFFFFF0;
    // rom_array[23787] = 32'hFFFFFFF0;
    // rom_array[23788] = 32'hFFFFFFF0;
    // rom_array[23789] = 32'hFFFFFFF1;
    // rom_array[23790] = 32'hFFFFFFF1;
    // rom_array[23791] = 32'hFFFFFFF1;
    // rom_array[23792] = 32'hFFFFFFF1;
    // rom_array[23793] = 32'hFFFFFFF0;
    // rom_array[23794] = 32'hFFFFFFF0;
    // rom_array[23795] = 32'hFFFFFFF0;
    // rom_array[23796] = 32'hFFFFFFF0;
    // rom_array[23797] = 32'hFFFFFFF1;
    // rom_array[23798] = 32'hFFFFFFF1;
    // rom_array[23799] = 32'hFFFFFFF1;
    // rom_array[23800] = 32'hFFFFFFF1;
    // rom_array[23801] = 32'hFFFFFFF0;
    // rom_array[23802] = 32'hFFFFFFF0;
    // rom_array[23803] = 32'hFFFFFFF0;
    // rom_array[23804] = 32'hFFFFFFF0;
    // rom_array[23805] = 32'hFFFFFFF1;
    // rom_array[23806] = 32'hFFFFFFF1;
    // rom_array[23807] = 32'hFFFFFFF1;
    // rom_array[23808] = 32'hFFFFFFF1;
    // rom_array[23809] = 32'hFFFFFFF0;
    // rom_array[23810] = 32'hFFFFFFF0;
    // rom_array[23811] = 32'hFFFFFFF0;
    // rom_array[23812] = 32'hFFFFFFF0;
    // rom_array[23813] = 32'hFFFFFFF1;
    // rom_array[23814] = 32'hFFFFFFF1;
    // rom_array[23815] = 32'hFFFFFFF1;
    // rom_array[23816] = 32'hFFFFFFF1;
    // rom_array[23817] = 32'hFFFFFFF0;
    // rom_array[23818] = 32'hFFFFFFF0;
    // rom_array[23819] = 32'hFFFFFFF0;
    // rom_array[23820] = 32'hFFFFFFF0;
    // rom_array[23821] = 32'hFFFFFFF1;
    // rom_array[23822] = 32'hFFFFFFF1;
    // rom_array[23823] = 32'hFFFFFFF1;
    // rom_array[23824] = 32'hFFFFFFF1;
    // rom_array[23825] = 32'hFFFFFFF0;
    // rom_array[23826] = 32'hFFFFFFF0;
    // rom_array[23827] = 32'hFFFFFFF0;
    // rom_array[23828] = 32'hFFFFFFF0;
    // rom_array[23829] = 32'hFFFFFFF1;
    // rom_array[23830] = 32'hFFFFFFF1;
    // rom_array[23831] = 32'hFFFFFFF1;
    // rom_array[23832] = 32'hFFFFFFF1;
    // rom_array[23833] = 32'hFFFFFFF1;
    // rom_array[23834] = 32'hFFFFFFF1;
    // rom_array[23835] = 32'hFFFFFFF1;
    // rom_array[23836] = 32'hFFFFFFF1;
    // rom_array[23837] = 32'hFFFFFFF1;
    // rom_array[23838] = 32'hFFFFFFF1;
    // rom_array[23839] = 32'hFFFFFFF1;
    // rom_array[23840] = 32'hFFFFFFF1;
    // rom_array[23841] = 32'hFFFFFFF1;
    // rom_array[23842] = 32'hFFFFFFF1;
    // rom_array[23843] = 32'hFFFFFFF1;
    // rom_array[23844] = 32'hFFFFFFF1;
    // rom_array[23845] = 32'hFFFFFFF1;
    // rom_array[23846] = 32'hFFFFFFF1;
    // rom_array[23847] = 32'hFFFFFFF1;
    // rom_array[23848] = 32'hFFFFFFF1;
    // rom_array[23849] = 32'hFFFFFFF1;
    // rom_array[23850] = 32'hFFFFFFF1;
    // rom_array[23851] = 32'hFFFFFFF1;
    // rom_array[23852] = 32'hFFFFFFF1;
    // rom_array[23853] = 32'hFFFFFFF1;
    // rom_array[23854] = 32'hFFFFFFF1;
    // rom_array[23855] = 32'hFFFFFFF1;
    // rom_array[23856] = 32'hFFFFFFF1;
    // rom_array[23857] = 32'hFFFFFFF1;
    // rom_array[23858] = 32'hFFFFFFF1;
    // rom_array[23859] = 32'hFFFFFFF1;
    // rom_array[23860] = 32'hFFFFFFF1;
    // rom_array[23861] = 32'hFFFFFFF1;
    // rom_array[23862] = 32'hFFFFFFF1;
    // rom_array[23863] = 32'hFFFFFFF1;
    // rom_array[23864] = 32'hFFFFFFF1;
    // rom_array[23865] = 32'hFFFFFFF1;
    // rom_array[23866] = 32'hFFFFFFF1;
    // rom_array[23867] = 32'hFFFFFFF1;
    // rom_array[23868] = 32'hFFFFFFF1;
    // rom_array[23869] = 32'hFFFFFFF1;
    // rom_array[23870] = 32'hFFFFFFF1;
    // rom_array[23871] = 32'hFFFFFFF1;
    // rom_array[23872] = 32'hFFFFFFF1;
    // rom_array[23873] = 32'hFFFFFFF1;
    // rom_array[23874] = 32'hFFFFFFF1;
    // rom_array[23875] = 32'hFFFFFFF1;
    // rom_array[23876] = 32'hFFFFFFF1;
    // rom_array[23877] = 32'hFFFFFFF1;
    // rom_array[23878] = 32'hFFFFFFF1;
    // rom_array[23879] = 32'hFFFFFFF1;
    // rom_array[23880] = 32'hFFFFFFF1;
    // rom_array[23881] = 32'hFFFFFFF1;
    // rom_array[23882] = 32'hFFFFFFF1;
    // rom_array[23883] = 32'hFFFFFFF1;
    // rom_array[23884] = 32'hFFFFFFF1;
    // rom_array[23885] = 32'hFFFFFFF1;
    // rom_array[23886] = 32'hFFFFFFF1;
    // rom_array[23887] = 32'hFFFFFFF1;
    // rom_array[23888] = 32'hFFFFFFF1;
    // rom_array[23889] = 32'hFFFFFFF1;
    // rom_array[23890] = 32'hFFFFFFF1;
    // rom_array[23891] = 32'hFFFFFFF1;
    // rom_array[23892] = 32'hFFFFFFF1;
    // rom_array[23893] = 32'hFFFFFFF1;
    // rom_array[23894] = 32'hFFFFFFF1;
    // rom_array[23895] = 32'hFFFFFFF1;
    // rom_array[23896] = 32'hFFFFFFF1;
    // rom_array[23897] = 32'hFFFFFFF1;
    // rom_array[23898] = 32'hFFFFFFF1;
    // rom_array[23899] = 32'hFFFFFFF1;
    // rom_array[23900] = 32'hFFFFFFF1;
    // rom_array[23901] = 32'hFFFFFFF1;
    // rom_array[23902] = 32'hFFFFFFF1;
    // rom_array[23903] = 32'hFFFFFFF1;
    // rom_array[23904] = 32'hFFFFFFF1;
    // rom_array[23905] = 32'hFFFFFFF1;
    // rom_array[23906] = 32'hFFFFFFF1;
    // rom_array[23907] = 32'hFFFFFFF1;
    // rom_array[23908] = 32'hFFFFFFF1;
    // rom_array[23909] = 32'hFFFFFFF1;
    // rom_array[23910] = 32'hFFFFFFF1;
    // rom_array[23911] = 32'hFFFFFFF1;
    // rom_array[23912] = 32'hFFFFFFF1;
    // rom_array[23913] = 32'hFFFFFFF1;
    // rom_array[23914] = 32'hFFFFFFF1;
    // rom_array[23915] = 32'hFFFFFFF1;
    // rom_array[23916] = 32'hFFFFFFF1;
    // rom_array[23917] = 32'hFFFFFFF1;
    // rom_array[23918] = 32'hFFFFFFF1;
    // rom_array[23919] = 32'hFFFFFFF1;
    // rom_array[23920] = 32'hFFFFFFF1;
    // rom_array[23921] = 32'hFFFFFFF1;
    // rom_array[23922] = 32'hFFFFFFF1;
    // rom_array[23923] = 32'hFFFFFFF1;
    // rom_array[23924] = 32'hFFFFFFF1;
    // rom_array[23925] = 32'hFFFFFFF1;
    // rom_array[23926] = 32'hFFFFFFF1;
    // rom_array[23927] = 32'hFFFFFFF1;
    // rom_array[23928] = 32'hFFFFFFF1;
    // rom_array[23929] = 32'hFFFFFFF1;
    // rom_array[23930] = 32'hFFFFFFF1;
    // rom_array[23931] = 32'hFFFFFFF1;
    // rom_array[23932] = 32'hFFFFFFF1;
    // rom_array[23933] = 32'hFFFFFFF1;
    // rom_array[23934] = 32'hFFFFFFF1;
    // rom_array[23935] = 32'hFFFFFFF1;
    // rom_array[23936] = 32'hFFFFFFF1;
    // rom_array[23937] = 32'hFFFFFFF1;
    // rom_array[23938] = 32'hFFFFFFF1;
    // rom_array[23939] = 32'hFFFFFFF1;
    // rom_array[23940] = 32'hFFFFFFF1;
    // rom_array[23941] = 32'hFFFFFFF1;
    // rom_array[23942] = 32'hFFFFFFF1;
    // rom_array[23943] = 32'hFFFFFFF1;
    // rom_array[23944] = 32'hFFFFFFF1;
    // rom_array[23945] = 32'hFFFFFFF1;
    // rom_array[23946] = 32'hFFFFFFF1;
    // rom_array[23947] = 32'hFFFFFFF1;
    // rom_array[23948] = 32'hFFFFFFF1;
    // rom_array[23949] = 32'hFFFFFFF1;
    // rom_array[23950] = 32'hFFFFFFF1;
    // rom_array[23951] = 32'hFFFFFFF1;
    // rom_array[23952] = 32'hFFFFFFF1;
    // rom_array[23953] = 32'hFFFFFFF1;
    // rom_array[23954] = 32'hFFFFFFF1;
    // rom_array[23955] = 32'hFFFFFFF1;
    // rom_array[23956] = 32'hFFFFFFF1;
    // rom_array[23957] = 32'hFFFFFFF1;
    // rom_array[23958] = 32'hFFFFFFF1;
    // rom_array[23959] = 32'hFFFFFFF1;
    // rom_array[23960] = 32'hFFFFFFF1;
    // rom_array[23961] = 32'hFFFFFFF1;
    // rom_array[23962] = 32'hFFFFFFF1;
    // rom_array[23963] = 32'hFFFFFFF1;
    // rom_array[23964] = 32'hFFFFFFF1;
    // rom_array[23965] = 32'hFFFFFFF1;
    // rom_array[23966] = 32'hFFFFFFF1;
    // rom_array[23967] = 32'hFFFFFFF1;
    // rom_array[23968] = 32'hFFFFFFF1;
    // rom_array[23969] = 32'hFFFFFFF1;
    // rom_array[23970] = 32'hFFFFFFF1;
    // rom_array[23971] = 32'hFFFFFFF1;
    // rom_array[23972] = 32'hFFFFFFF1;
    // rom_array[23973] = 32'hFFFFFFF1;
    // rom_array[23974] = 32'hFFFFFFF1;
    // rom_array[23975] = 32'hFFFFFFF1;
    // rom_array[23976] = 32'hFFFFFFF1;
    // rom_array[23977] = 32'hFFFFFFF1;
    // rom_array[23978] = 32'hFFFFFFF1;
    // rom_array[23979] = 32'hFFFFFFF1;
    // rom_array[23980] = 32'hFFFFFFF1;
    // rom_array[23981] = 32'hFFFFFFF1;
    // rom_array[23982] = 32'hFFFFFFF1;
    // rom_array[23983] = 32'hFFFFFFF1;
    // rom_array[23984] = 32'hFFFFFFF1;
    // rom_array[23985] = 32'hFFFFFFF1;
    // rom_array[23986] = 32'hFFFFFFF1;
    // rom_array[23987] = 32'hFFFFFFF1;
    // rom_array[23988] = 32'hFFFFFFF1;
    // rom_array[23989] = 32'hFFFFFFF1;
    // rom_array[23990] = 32'hFFFFFFF1;
    // rom_array[23991] = 32'hFFFFFFF1;
    // rom_array[23992] = 32'hFFFFFFF1;
    // rom_array[23993] = 32'hFFFFFFF1;
    // rom_array[23994] = 32'hFFFFFFF1;
    // rom_array[23995] = 32'hFFFFFFF1;
    // rom_array[23996] = 32'hFFFFFFF1;
    // rom_array[23997] = 32'hFFFFFFF1;
    // rom_array[23998] = 32'hFFFFFFF1;
    // rom_array[23999] = 32'hFFFFFFF1;
    // rom_array[24000] = 32'hFFFFFFF1;
    // rom_array[24001] = 32'hFFFFFFF1;
    // rom_array[24002] = 32'hFFFFFFF1;
    // rom_array[24003] = 32'hFFFFFFF1;
    // rom_array[24004] = 32'hFFFFFFF1;
    // rom_array[24005] = 32'hFFFFFFF1;
    // rom_array[24006] = 32'hFFFFFFF1;
    // rom_array[24007] = 32'hFFFFFFF1;
    // rom_array[24008] = 32'hFFFFFFF1;
    // rom_array[24009] = 32'hFFFFFFF1;
    // rom_array[24010] = 32'hFFFFFFF1;
    // rom_array[24011] = 32'hFFFFFFF1;
    // rom_array[24012] = 32'hFFFFFFF1;
    // rom_array[24013] = 32'hFFFFFFF1;
    // rom_array[24014] = 32'hFFFFFFF1;
    // rom_array[24015] = 32'hFFFFFFF1;
    // rom_array[24016] = 32'hFFFFFFF1;
    // rom_array[24017] = 32'hFFFFFFF1;
    // rom_array[24018] = 32'hFFFFFFF1;
    // rom_array[24019] = 32'hFFFFFFF1;
    // rom_array[24020] = 32'hFFFFFFF1;
    // rom_array[24021] = 32'hFFFFFFF1;
    // rom_array[24022] = 32'hFFFFFFF1;
    // rom_array[24023] = 32'hFFFFFFF1;
    // rom_array[24024] = 32'hFFFFFFF1;
    // rom_array[24025] = 32'hFFFFFFF1;
    // rom_array[24026] = 32'hFFFFFFF1;
    // rom_array[24027] = 32'hFFFFFFF1;
    // rom_array[24028] = 32'hFFFFFFF1;
    // rom_array[24029] = 32'hFFFFFFF1;
    // rom_array[24030] = 32'hFFFFFFF1;
    // rom_array[24031] = 32'hFFFFFFF1;
    // rom_array[24032] = 32'hFFFFFFF1;
    // rom_array[24033] = 32'hFFFFFFF1;
    // rom_array[24034] = 32'hFFFFFFF1;
    // rom_array[24035] = 32'hFFFFFFF1;
    // rom_array[24036] = 32'hFFFFFFF1;
    // rom_array[24037] = 32'hFFFFFFF1;
    // rom_array[24038] = 32'hFFFFFFF1;
    // rom_array[24039] = 32'hFFFFFFF1;
    // rom_array[24040] = 32'hFFFFFFF1;
    // rom_array[24041] = 32'hFFFFFFF0;
    // rom_array[24042] = 32'hFFFFFFF0;
    // rom_array[24043] = 32'hFFFFFFF0;
    // rom_array[24044] = 32'hFFFFFFF0;
    // rom_array[24045] = 32'hFFFFFFF1;
    // rom_array[24046] = 32'hFFFFFFF1;
    // rom_array[24047] = 32'hFFFFFFF1;
    // rom_array[24048] = 32'hFFFFFFF1;
    // rom_array[24049] = 32'hFFFFFFF0;
    // rom_array[24050] = 32'hFFFFFFF0;
    // rom_array[24051] = 32'hFFFFFFF0;
    // rom_array[24052] = 32'hFFFFFFF0;
    // rom_array[24053] = 32'hFFFFFFF1;
    // rom_array[24054] = 32'hFFFFFFF1;
    // rom_array[24055] = 32'hFFFFFFF1;
    // rom_array[24056] = 32'hFFFFFFF1;
    // rom_array[24057] = 32'hFFFFFFF0;
    // rom_array[24058] = 32'hFFFFFFF0;
    // rom_array[24059] = 32'hFFFFFFF0;
    // rom_array[24060] = 32'hFFFFFFF0;
    // rom_array[24061] = 32'hFFFFFFF1;
    // rom_array[24062] = 32'hFFFFFFF1;
    // rom_array[24063] = 32'hFFFFFFF1;
    // rom_array[24064] = 32'hFFFFFFF1;
    // rom_array[24065] = 32'hFFFFFFF0;
    // rom_array[24066] = 32'hFFFFFFF0;
    // rom_array[24067] = 32'hFFFFFFF0;
    // rom_array[24068] = 32'hFFFFFFF0;
    // rom_array[24069] = 32'hFFFFFFF1;
    // rom_array[24070] = 32'hFFFFFFF1;
    // rom_array[24071] = 32'hFFFFFFF1;
    // rom_array[24072] = 32'hFFFFFFF1;
    // rom_array[24073] = 32'hFFFFFFF0;
    // rom_array[24074] = 32'hFFFFFFF0;
    // rom_array[24075] = 32'hFFFFFFF0;
    // rom_array[24076] = 32'hFFFFFFF0;
    // rom_array[24077] = 32'hFFFFFFF1;
    // rom_array[24078] = 32'hFFFFFFF1;
    // rom_array[24079] = 32'hFFFFFFF1;
    // rom_array[24080] = 32'hFFFFFFF1;
    // rom_array[24081] = 32'hFFFFFFF0;
    // rom_array[24082] = 32'hFFFFFFF0;
    // rom_array[24083] = 32'hFFFFFFF0;
    // rom_array[24084] = 32'hFFFFFFF0;
    // rom_array[24085] = 32'hFFFFFFF1;
    // rom_array[24086] = 32'hFFFFFFF1;
    // rom_array[24087] = 32'hFFFFFFF1;
    // rom_array[24088] = 32'hFFFFFFF1;
    // rom_array[24089] = 32'hFFFFFFF0;
    // rom_array[24090] = 32'hFFFFFFF0;
    // rom_array[24091] = 32'hFFFFFFF1;
    // rom_array[24092] = 32'hFFFFFFF1;
    // rom_array[24093] = 32'hFFFFFFF0;
    // rom_array[24094] = 32'hFFFFFFF0;
    // rom_array[24095] = 32'hFFFFFFF1;
    // rom_array[24096] = 32'hFFFFFFF1;
    // rom_array[24097] = 32'hFFFFFFF0;
    // rom_array[24098] = 32'hFFFFFFF0;
    // rom_array[24099] = 32'hFFFFFFF1;
    // rom_array[24100] = 32'hFFFFFFF1;
    // rom_array[24101] = 32'hFFFFFFF0;
    // rom_array[24102] = 32'hFFFFFFF0;
    // rom_array[24103] = 32'hFFFFFFF1;
    // rom_array[24104] = 32'hFFFFFFF1;
    // rom_array[24105] = 32'hFFFFFFF0;
    // rom_array[24106] = 32'hFFFFFFF0;
    // rom_array[24107] = 32'hFFFFFFF1;
    // rom_array[24108] = 32'hFFFFFFF1;
    // rom_array[24109] = 32'hFFFFFFF0;
    // rom_array[24110] = 32'hFFFFFFF0;
    // rom_array[24111] = 32'hFFFFFFF1;
    // rom_array[24112] = 32'hFFFFFFF1;
    // rom_array[24113] = 32'hFFFFFFF0;
    // rom_array[24114] = 32'hFFFFFFF0;
    // rom_array[24115] = 32'hFFFFFFF1;
    // rom_array[24116] = 32'hFFFFFFF1;
    // rom_array[24117] = 32'hFFFFFFF0;
    // rom_array[24118] = 32'hFFFFFFF0;
    // rom_array[24119] = 32'hFFFFFFF1;
    // rom_array[24120] = 32'hFFFFFFF1;
    // rom_array[24121] = 32'hFFFFFFF0;
    // rom_array[24122] = 32'hFFFFFFF0;
    // rom_array[24123] = 32'hFFFFFFF0;
    // rom_array[24124] = 32'hFFFFFFF0;
    // rom_array[24125] = 32'hFFFFFFF1;
    // rom_array[24126] = 32'hFFFFFFF1;
    // rom_array[24127] = 32'hFFFFFFF1;
    // rom_array[24128] = 32'hFFFFFFF1;
    // rom_array[24129] = 32'hFFFFFFF0;
    // rom_array[24130] = 32'hFFFFFFF0;
    // rom_array[24131] = 32'hFFFFFFF0;
    // rom_array[24132] = 32'hFFFFFFF0;
    // rom_array[24133] = 32'hFFFFFFF1;
    // rom_array[24134] = 32'hFFFFFFF1;
    // rom_array[24135] = 32'hFFFFFFF1;
    // rom_array[24136] = 32'hFFFFFFF1;
    // rom_array[24137] = 32'hFFFFFFF0;
    // rom_array[24138] = 32'hFFFFFFF0;
    // rom_array[24139] = 32'hFFFFFFF0;
    // rom_array[24140] = 32'hFFFFFFF0;
    // rom_array[24141] = 32'hFFFFFFF1;
    // rom_array[24142] = 32'hFFFFFFF1;
    // rom_array[24143] = 32'hFFFFFFF1;
    // rom_array[24144] = 32'hFFFFFFF1;
    // rom_array[24145] = 32'hFFFFFFF0;
    // rom_array[24146] = 32'hFFFFFFF0;
    // rom_array[24147] = 32'hFFFFFFF0;
    // rom_array[24148] = 32'hFFFFFFF0;
    // rom_array[24149] = 32'hFFFFFFF1;
    // rom_array[24150] = 32'hFFFFFFF1;
    // rom_array[24151] = 32'hFFFFFFF1;
    // rom_array[24152] = 32'hFFFFFFF1;
    // rom_array[24153] = 32'hFFFFFFF0;
    // rom_array[24154] = 32'hFFFFFFF0;
    // rom_array[24155] = 32'hFFFFFFF1;
    // rom_array[24156] = 32'hFFFFFFF1;
    // rom_array[24157] = 32'hFFFFFFF0;
    // rom_array[24158] = 32'hFFFFFFF0;
    // rom_array[24159] = 32'hFFFFFFF1;
    // rom_array[24160] = 32'hFFFFFFF1;
    // rom_array[24161] = 32'hFFFFFFF0;
    // rom_array[24162] = 32'hFFFFFFF0;
    // rom_array[24163] = 32'hFFFFFFF1;
    // rom_array[24164] = 32'hFFFFFFF1;
    // rom_array[24165] = 32'hFFFFFFF0;
    // rom_array[24166] = 32'hFFFFFFF0;
    // rom_array[24167] = 32'hFFFFFFF1;
    // rom_array[24168] = 32'hFFFFFFF1;
    // rom_array[24169] = 32'hFFFFFFF0;
    // rom_array[24170] = 32'hFFFFFFF0;
    // rom_array[24171] = 32'hFFFFFFF1;
    // rom_array[24172] = 32'hFFFFFFF1;
    // rom_array[24173] = 32'hFFFFFFF1;
    // rom_array[24174] = 32'hFFFFFFF1;
    // rom_array[24175] = 32'hFFFFFFF1;
    // rom_array[24176] = 32'hFFFFFFF1;
    // rom_array[24177] = 32'hFFFFFFF0;
    // rom_array[24178] = 32'hFFFFFFF0;
    // rom_array[24179] = 32'hFFFFFFF1;
    // rom_array[24180] = 32'hFFFFFFF1;
    // rom_array[24181] = 32'hFFFFFFF1;
    // rom_array[24182] = 32'hFFFFFFF1;
    // rom_array[24183] = 32'hFFFFFFF1;
    // rom_array[24184] = 32'hFFFFFFF1;
    // rom_array[24185] = 32'hFFFFFFF0;
    // rom_array[24186] = 32'hFFFFFFF0;
    // rom_array[24187] = 32'hFFFFFFF0;
    // rom_array[24188] = 32'hFFFFFFF0;
    // rom_array[24189] = 32'hFFFFFFF1;
    // rom_array[24190] = 32'hFFFFFFF1;
    // rom_array[24191] = 32'hFFFFFFF1;
    // rom_array[24192] = 32'hFFFFFFF1;
    // rom_array[24193] = 32'hFFFFFFF0;
    // rom_array[24194] = 32'hFFFFFFF0;
    // rom_array[24195] = 32'hFFFFFFF0;
    // rom_array[24196] = 32'hFFFFFFF0;
    // rom_array[24197] = 32'hFFFFFFF1;
    // rom_array[24198] = 32'hFFFFFFF1;
    // rom_array[24199] = 32'hFFFFFFF1;
    // rom_array[24200] = 32'hFFFFFFF1;
    // rom_array[24201] = 32'hFFFFFFF1;
    // rom_array[24202] = 32'hFFFFFFF1;
    // rom_array[24203] = 32'hFFFFFFF1;
    // rom_array[24204] = 32'hFFFFFFF1;
    // rom_array[24205] = 32'hFFFFFFF0;
    // rom_array[24206] = 32'hFFFFFFF0;
    // rom_array[24207] = 32'hFFFFFFF0;
    // rom_array[24208] = 32'hFFFFFFF0;
    // rom_array[24209] = 32'hFFFFFFF1;
    // rom_array[24210] = 32'hFFFFFFF1;
    // rom_array[24211] = 32'hFFFFFFF1;
    // rom_array[24212] = 32'hFFFFFFF1;
    // rom_array[24213] = 32'hFFFFFFF0;
    // rom_array[24214] = 32'hFFFFFFF0;
    // rom_array[24215] = 32'hFFFFFFF0;
    // rom_array[24216] = 32'hFFFFFFF0;
    // rom_array[24217] = 32'hFFFFFFF1;
    // rom_array[24218] = 32'hFFFFFFF1;
    // rom_array[24219] = 32'hFFFFFFF1;
    // rom_array[24220] = 32'hFFFFFFF1;
    // rom_array[24221] = 32'hFFFFFFF0;
    // rom_array[24222] = 32'hFFFFFFF0;
    // rom_array[24223] = 32'hFFFFFFF0;
    // rom_array[24224] = 32'hFFFFFFF0;
    // rom_array[24225] = 32'hFFFFFFF1;
    // rom_array[24226] = 32'hFFFFFFF1;
    // rom_array[24227] = 32'hFFFFFFF1;
    // rom_array[24228] = 32'hFFFFFFF1;
    // rom_array[24229] = 32'hFFFFFFF0;
    // rom_array[24230] = 32'hFFFFFFF0;
    // rom_array[24231] = 32'hFFFFFFF0;
    // rom_array[24232] = 32'hFFFFFFF0;
    // rom_array[24233] = 32'hFFFFFFF1;
    // rom_array[24234] = 32'hFFFFFFF1;
    // rom_array[24235] = 32'hFFFFFFF1;
    // rom_array[24236] = 32'hFFFFFFF1;
    // rom_array[24237] = 32'hFFFFFFF0;
    // rom_array[24238] = 32'hFFFFFFF0;
    // rom_array[24239] = 32'hFFFFFFF0;
    // rom_array[24240] = 32'hFFFFFFF0;
    // rom_array[24241] = 32'hFFFFFFF1;
    // rom_array[24242] = 32'hFFFFFFF1;
    // rom_array[24243] = 32'hFFFFFFF1;
    // rom_array[24244] = 32'hFFFFFFF1;
    // rom_array[24245] = 32'hFFFFFFF0;
    // rom_array[24246] = 32'hFFFFFFF0;
    // rom_array[24247] = 32'hFFFFFFF0;
    // rom_array[24248] = 32'hFFFFFFF0;
    // rom_array[24249] = 32'hFFFFFFF1;
    // rom_array[24250] = 32'hFFFFFFF1;
    // rom_array[24251] = 32'hFFFFFFF1;
    // rom_array[24252] = 32'hFFFFFFF1;
    // rom_array[24253] = 32'hFFFFFFF0;
    // rom_array[24254] = 32'hFFFFFFF0;
    // rom_array[24255] = 32'hFFFFFFF0;
    // rom_array[24256] = 32'hFFFFFFF0;
    // rom_array[24257] = 32'hFFFFFFF1;
    // rom_array[24258] = 32'hFFFFFFF1;
    // rom_array[24259] = 32'hFFFFFFF1;
    // rom_array[24260] = 32'hFFFFFFF1;
    // rom_array[24261] = 32'hFFFFFFF0;
    // rom_array[24262] = 32'hFFFFFFF0;
    // rom_array[24263] = 32'hFFFFFFF0;
    // rom_array[24264] = 32'hFFFFFFF0;
    // rom_array[24265] = 32'hFFFFFFF1;
    // rom_array[24266] = 32'hFFFFFFF1;
    // rom_array[24267] = 32'hFFFFFFF1;
    // rom_array[24268] = 32'hFFFFFFF1;
    // rom_array[24269] = 32'hFFFFFFF0;
    // rom_array[24270] = 32'hFFFFFFF0;
    // rom_array[24271] = 32'hFFFFFFF0;
    // rom_array[24272] = 32'hFFFFFFF0;
    // rom_array[24273] = 32'hFFFFFFF1;
    // rom_array[24274] = 32'hFFFFFFF1;
    // rom_array[24275] = 32'hFFFFFFF1;
    // rom_array[24276] = 32'hFFFFFFF1;
    // rom_array[24277] = 32'hFFFFFFF0;
    // rom_array[24278] = 32'hFFFFFFF0;
    // rom_array[24279] = 32'hFFFFFFF0;
    // rom_array[24280] = 32'hFFFFFFF0;
    // rom_array[24281] = 32'hFFFFFFF0;
    // rom_array[24282] = 32'hFFFFFFF0;
    // rom_array[24283] = 32'hFFFFFFF1;
    // rom_array[24284] = 32'hFFFFFFF1;
    // rom_array[24285] = 32'hFFFFFFF0;
    // rom_array[24286] = 32'hFFFFFFF0;
    // rom_array[24287] = 32'hFFFFFFF0;
    // rom_array[24288] = 32'hFFFFFFF0;
    // rom_array[24289] = 32'hFFFFFFF0;
    // rom_array[24290] = 32'hFFFFFFF0;
    // rom_array[24291] = 32'hFFFFFFF1;
    // rom_array[24292] = 32'hFFFFFFF1;
    // rom_array[24293] = 32'hFFFFFFF0;
    // rom_array[24294] = 32'hFFFFFFF0;
    // rom_array[24295] = 32'hFFFFFFF0;
    // rom_array[24296] = 32'hFFFFFFF0;
    // rom_array[24297] = 32'hFFFFFFF1;
    // rom_array[24298] = 32'hFFFFFFF1;
    // rom_array[24299] = 32'hFFFFFFF1;
    // rom_array[24300] = 32'hFFFFFFF1;
    // rom_array[24301] = 32'hFFFFFFF1;
    // rom_array[24302] = 32'hFFFFFFF1;
    // rom_array[24303] = 32'hFFFFFFF1;
    // rom_array[24304] = 32'hFFFFFFF1;
    // rom_array[24305] = 32'hFFFFFFF1;
    // rom_array[24306] = 32'hFFFFFFF1;
    // rom_array[24307] = 32'hFFFFFFF1;
    // rom_array[24308] = 32'hFFFFFFF1;
    // rom_array[24309] = 32'hFFFFFFF1;
    // rom_array[24310] = 32'hFFFFFFF1;
    // rom_array[24311] = 32'hFFFFFFF1;
    // rom_array[24312] = 32'hFFFFFFF1;
    // rom_array[24313] = 32'hFFFFFFF1;
    // rom_array[24314] = 32'hFFFFFFF1;
    // rom_array[24315] = 32'hFFFFFFF1;
    // rom_array[24316] = 32'hFFFFFFF1;
    // rom_array[24317] = 32'hFFFFFFF1;
    // rom_array[24318] = 32'hFFFFFFF1;
    // rom_array[24319] = 32'hFFFFFFF1;
    // rom_array[24320] = 32'hFFFFFFF1;
    // rom_array[24321] = 32'hFFFFFFF1;
    // rom_array[24322] = 32'hFFFFFFF1;
    // rom_array[24323] = 32'hFFFFFFF1;
    // rom_array[24324] = 32'hFFFFFFF1;
    // rom_array[24325] = 32'hFFFFFFF1;
    // rom_array[24326] = 32'hFFFFFFF1;
    // rom_array[24327] = 32'hFFFFFFF1;
    // rom_array[24328] = 32'hFFFFFFF1;
    // rom_array[24329] = 32'hFFFFFFF1;
    // rom_array[24330] = 32'hFFFFFFF1;
    // rom_array[24331] = 32'hFFFFFFF1;
    // rom_array[24332] = 32'hFFFFFFF1;
    // rom_array[24333] = 32'hFFFFFFF0;
    // rom_array[24334] = 32'hFFFFFFF0;
    // rom_array[24335] = 32'hFFFFFFF0;
    // rom_array[24336] = 32'hFFFFFFF0;
    // rom_array[24337] = 32'hFFFFFFF1;
    // rom_array[24338] = 32'hFFFFFFF1;
    // rom_array[24339] = 32'hFFFFFFF1;
    // rom_array[24340] = 32'hFFFFFFF1;
    // rom_array[24341] = 32'hFFFFFFF0;
    // rom_array[24342] = 32'hFFFFFFF0;
    // rom_array[24343] = 32'hFFFFFFF0;
    // rom_array[24344] = 32'hFFFFFFF0;
    // rom_array[24345] = 32'hFFFFFFF1;
    // rom_array[24346] = 32'hFFFFFFF1;
    // rom_array[24347] = 32'hFFFFFFF1;
    // rom_array[24348] = 32'hFFFFFFF1;
    // rom_array[24349] = 32'hFFFFFFF0;
    // rom_array[24350] = 32'hFFFFFFF0;
    // rom_array[24351] = 32'hFFFFFFF0;
    // rom_array[24352] = 32'hFFFFFFF0;
    // rom_array[24353] = 32'hFFFFFFF1;
    // rom_array[24354] = 32'hFFFFFFF1;
    // rom_array[24355] = 32'hFFFFFFF1;
    // rom_array[24356] = 32'hFFFFFFF1;
    // rom_array[24357] = 32'hFFFFFFF0;
    // rom_array[24358] = 32'hFFFFFFF0;
    // rom_array[24359] = 32'hFFFFFFF0;
    // rom_array[24360] = 32'hFFFFFFF0;
    // rom_array[24361] = 32'hFFFFFFF1;
    // rom_array[24362] = 32'hFFFFFFF1;
    // rom_array[24363] = 32'hFFFFFFF1;
    // rom_array[24364] = 32'hFFFFFFF1;
    // rom_array[24365] = 32'hFFFFFFF1;
    // rom_array[24366] = 32'hFFFFFFF1;
    // rom_array[24367] = 32'hFFFFFFF1;
    // rom_array[24368] = 32'hFFFFFFF1;
    // rom_array[24369] = 32'hFFFFFFF1;
    // rom_array[24370] = 32'hFFFFFFF1;
    // rom_array[24371] = 32'hFFFFFFF1;
    // rom_array[24372] = 32'hFFFFFFF1;
    // rom_array[24373] = 32'hFFFFFFF1;
    // rom_array[24374] = 32'hFFFFFFF1;
    // rom_array[24375] = 32'hFFFFFFF1;
    // rom_array[24376] = 32'hFFFFFFF1;
    // rom_array[24377] = 32'hFFFFFFF1;
    // rom_array[24378] = 32'hFFFFFFF1;
    // rom_array[24379] = 32'hFFFFFFF1;
    // rom_array[24380] = 32'hFFFFFFF1;
    // rom_array[24381] = 32'hFFFFFFF0;
    // rom_array[24382] = 32'hFFFFFFF0;
    // rom_array[24383] = 32'hFFFFFFF0;
    // rom_array[24384] = 32'hFFFFFFF0;
    // rom_array[24385] = 32'hFFFFFFF1;
    // rom_array[24386] = 32'hFFFFFFF1;
    // rom_array[24387] = 32'hFFFFFFF1;
    // rom_array[24388] = 32'hFFFFFFF1;
    // rom_array[24389] = 32'hFFFFFFF0;
    // rom_array[24390] = 32'hFFFFFFF0;
    // rom_array[24391] = 32'hFFFFFFF0;
    // rom_array[24392] = 32'hFFFFFFF0;
    // rom_array[24393] = 32'hFFFFFFF1;
    // rom_array[24394] = 32'hFFFFFFF1;
    // rom_array[24395] = 32'hFFFFFFF1;
    // rom_array[24396] = 32'hFFFFFFF1;
    // rom_array[24397] = 32'hFFFFFFF0;
    // rom_array[24398] = 32'hFFFFFFF0;
    // rom_array[24399] = 32'hFFFFFFF0;
    // rom_array[24400] = 32'hFFFFFFF0;
    // rom_array[24401] = 32'hFFFFFFF1;
    // rom_array[24402] = 32'hFFFFFFF1;
    // rom_array[24403] = 32'hFFFFFFF1;
    // rom_array[24404] = 32'hFFFFFFF1;
    // rom_array[24405] = 32'hFFFFFFF0;
    // rom_array[24406] = 32'hFFFFFFF0;
    // rom_array[24407] = 32'hFFFFFFF0;
    // rom_array[24408] = 32'hFFFFFFF0;
    // rom_array[24409] = 32'hFFFFFFF1;
    // rom_array[24410] = 32'hFFFFFFF1;
    // rom_array[24411] = 32'hFFFFFFF1;
    // rom_array[24412] = 32'hFFFFFFF1;
    // rom_array[24413] = 32'hFFFFFFF1;
    // rom_array[24414] = 32'hFFFFFFF1;
    // rom_array[24415] = 32'hFFFFFFF1;
    // rom_array[24416] = 32'hFFFFFFF1;
    // rom_array[24417] = 32'hFFFFFFF1;
    // rom_array[24418] = 32'hFFFFFFF1;
    // rom_array[24419] = 32'hFFFFFFF1;
    // rom_array[24420] = 32'hFFFFFFF1;
    // rom_array[24421] = 32'hFFFFFFF1;
    // rom_array[24422] = 32'hFFFFFFF1;
    // rom_array[24423] = 32'hFFFFFFF1;
    // rom_array[24424] = 32'hFFFFFFF1;
    // rom_array[24425] = 32'hFFFFFFF1;
    // rom_array[24426] = 32'hFFFFFFF1;
    // rom_array[24427] = 32'hFFFFFFF1;
    // rom_array[24428] = 32'hFFFFFFF1;
    // rom_array[24429] = 32'hFFFFFFF1;
    // rom_array[24430] = 32'hFFFFFFF1;
    // rom_array[24431] = 32'hFFFFFFF1;
    // rom_array[24432] = 32'hFFFFFFF1;
    // rom_array[24433] = 32'hFFFFFFF1;
    // rom_array[24434] = 32'hFFFFFFF1;
    // rom_array[24435] = 32'hFFFFFFF1;
    // rom_array[24436] = 32'hFFFFFFF1;
    // rom_array[24437] = 32'hFFFFFFF1;
    // rom_array[24438] = 32'hFFFFFFF1;
    // rom_array[24439] = 32'hFFFFFFF1;
    // rom_array[24440] = 32'hFFFFFFF1;
    // rom_array[24441] = 32'hFFFFFFF1;
    // rom_array[24442] = 32'hFFFFFFF1;
    // rom_array[24443] = 32'hFFFFFFF1;
    // rom_array[24444] = 32'hFFFFFFF1;
    // rom_array[24445] = 32'hFFFFFFF1;
    // rom_array[24446] = 32'hFFFFFFF1;
    // rom_array[24447] = 32'hFFFFFFF1;
    // rom_array[24448] = 32'hFFFFFFF1;
    // rom_array[24449] = 32'hFFFFFFF1;
    // rom_array[24450] = 32'hFFFFFFF1;
    // rom_array[24451] = 32'hFFFFFFF1;
    // rom_array[24452] = 32'hFFFFFFF1;
    // rom_array[24453] = 32'hFFFFFFF1;
    // rom_array[24454] = 32'hFFFFFFF1;
    // rom_array[24455] = 32'hFFFFFFF1;
    // rom_array[24456] = 32'hFFFFFFF1;
    // rom_array[24457] = 32'hFFFFFFF1;
    // rom_array[24458] = 32'hFFFFFFF1;
    // rom_array[24459] = 32'hFFFFFFF1;
    // rom_array[24460] = 32'hFFFFFFF1;
    // rom_array[24461] = 32'hFFFFFFF1;
    // rom_array[24462] = 32'hFFFFFFF1;
    // rom_array[24463] = 32'hFFFFFFF1;
    // rom_array[24464] = 32'hFFFFFFF1;
    // rom_array[24465] = 32'hFFFFFFF1;
    // rom_array[24466] = 32'hFFFFFFF1;
    // rom_array[24467] = 32'hFFFFFFF1;
    // rom_array[24468] = 32'hFFFFFFF1;
    // rom_array[24469] = 32'hFFFFFFF1;
    // rom_array[24470] = 32'hFFFFFFF1;
    // rom_array[24471] = 32'hFFFFFFF1;
    // rom_array[24472] = 32'hFFFFFFF1;
    // rom_array[24473] = 32'hFFFFFFF1;
    // rom_array[24474] = 32'hFFFFFFF1;
    // rom_array[24475] = 32'hFFFFFFF1;
    // rom_array[24476] = 32'hFFFFFFF1;
    // rom_array[24477] = 32'hFFFFFFF0;
    // rom_array[24478] = 32'hFFFFFFF0;
    // rom_array[24479] = 32'hFFFFFFF0;
    // rom_array[24480] = 32'hFFFFFFF0;
    // rom_array[24481] = 32'hFFFFFFF1;
    // rom_array[24482] = 32'hFFFFFFF1;
    // rom_array[24483] = 32'hFFFFFFF1;
    // rom_array[24484] = 32'hFFFFFFF1;
    // rom_array[24485] = 32'hFFFFFFF0;
    // rom_array[24486] = 32'hFFFFFFF0;
    // rom_array[24487] = 32'hFFFFFFF0;
    // rom_array[24488] = 32'hFFFFFFF0;
    // rom_array[24489] = 32'hFFFFFFF1;
    // rom_array[24490] = 32'hFFFFFFF1;
    // rom_array[24491] = 32'hFFFFFFF1;
    // rom_array[24492] = 32'hFFFFFFF1;
    // rom_array[24493] = 32'hFFFFFFF0;
    // rom_array[24494] = 32'hFFFFFFF0;
    // rom_array[24495] = 32'hFFFFFFF0;
    // rom_array[24496] = 32'hFFFFFFF0;
    // rom_array[24497] = 32'hFFFFFFF1;
    // rom_array[24498] = 32'hFFFFFFF1;
    // rom_array[24499] = 32'hFFFFFFF1;
    // rom_array[24500] = 32'hFFFFFFF1;
    // rom_array[24501] = 32'hFFFFFFF0;
    // rom_array[24502] = 32'hFFFFFFF0;
    // rom_array[24503] = 32'hFFFFFFF0;
    // rom_array[24504] = 32'hFFFFFFF0;
    // rom_array[24505] = 32'hFFFFFFF1;
    // rom_array[24506] = 32'hFFFFFFF1;
    // rom_array[24507] = 32'hFFFFFFF1;
    // rom_array[24508] = 32'hFFFFFFF1;
    // rom_array[24509] = 32'hFFFFFFF0;
    // rom_array[24510] = 32'hFFFFFFF0;
    // rom_array[24511] = 32'hFFFFFFF0;
    // rom_array[24512] = 32'hFFFFFFF0;
    // rom_array[24513] = 32'hFFFFFFF1;
    // rom_array[24514] = 32'hFFFFFFF1;
    // rom_array[24515] = 32'hFFFFFFF1;
    // rom_array[24516] = 32'hFFFFFFF1;
    // rom_array[24517] = 32'hFFFFFFF0;
    // rom_array[24518] = 32'hFFFFFFF0;
    // rom_array[24519] = 32'hFFFFFFF0;
    // rom_array[24520] = 32'hFFFFFFF0;
    // rom_array[24521] = 32'hFFFFFFF0;
    // rom_array[24522] = 32'hFFFFFFF0;
    // rom_array[24523] = 32'hFFFFFFF0;
    // rom_array[24524] = 32'hFFFFFFF0;
    // rom_array[24525] = 32'hFFFFFFF1;
    // rom_array[24526] = 32'hFFFFFFF1;
    // rom_array[24527] = 32'hFFFFFFF1;
    // rom_array[24528] = 32'hFFFFFFF1;
    // rom_array[24529] = 32'hFFFFFFF0;
    // rom_array[24530] = 32'hFFFFFFF0;
    // rom_array[24531] = 32'hFFFFFFF0;
    // rom_array[24532] = 32'hFFFFFFF0;
    // rom_array[24533] = 32'hFFFFFFF1;
    // rom_array[24534] = 32'hFFFFFFF1;
    // rom_array[24535] = 32'hFFFFFFF1;
    // rom_array[24536] = 32'hFFFFFFF1;
    // rom_array[24537] = 32'hFFFFFFF0;
    // rom_array[24538] = 32'hFFFFFFF0;
    // rom_array[24539] = 32'hFFFFFFF0;
    // rom_array[24540] = 32'hFFFFFFF0;
    // rom_array[24541] = 32'hFFFFFFF1;
    // rom_array[24542] = 32'hFFFFFFF1;
    // rom_array[24543] = 32'hFFFFFFF1;
    // rom_array[24544] = 32'hFFFFFFF1;
    // rom_array[24545] = 32'hFFFFFFF0;
    // rom_array[24546] = 32'hFFFFFFF0;
    // rom_array[24547] = 32'hFFFFFFF0;
    // rom_array[24548] = 32'hFFFFFFF0;
    // rom_array[24549] = 32'hFFFFFFF1;
    // rom_array[24550] = 32'hFFFFFFF1;
    // rom_array[24551] = 32'hFFFFFFF1;
    // rom_array[24552] = 32'hFFFFFFF1;
    // rom_array[24553] = 32'hFFFFFFF0;
    // rom_array[24554] = 32'hFFFFFFF0;
    // rom_array[24555] = 32'hFFFFFFF0;
    // rom_array[24556] = 32'hFFFFFFF0;
    // rom_array[24557] = 32'hFFFFFFF1;
    // rom_array[24558] = 32'hFFFFFFF1;
    // rom_array[24559] = 32'hFFFFFFF1;
    // rom_array[24560] = 32'hFFFFFFF1;
    // rom_array[24561] = 32'hFFFFFFF0;
    // rom_array[24562] = 32'hFFFFFFF0;
    // rom_array[24563] = 32'hFFFFFFF0;
    // rom_array[24564] = 32'hFFFFFFF0;
    // rom_array[24565] = 32'hFFFFFFF1;
    // rom_array[24566] = 32'hFFFFFFF1;
    // rom_array[24567] = 32'hFFFFFFF1;
    // rom_array[24568] = 32'hFFFFFFF1;
    // rom_array[24569] = 32'hFFFFFFF0;
    // rom_array[24570] = 32'hFFFFFFF0;
    // rom_array[24571] = 32'hFFFFFFF0;
    // rom_array[24572] = 32'hFFFFFFF0;
    // rom_array[24573] = 32'hFFFFFFF1;
    // rom_array[24574] = 32'hFFFFFFF1;
    // rom_array[24575] = 32'hFFFFFFF1;
    // rom_array[24576] = 32'hFFFFFFF1;
    // rom_array[24577] = 32'hFFFFFFF0;
    // rom_array[24578] = 32'hFFFFFFF0;
    // rom_array[24579] = 32'hFFFFFFF0;
    // rom_array[24580] = 32'hFFFFFFF0;
    // rom_array[24581] = 32'hFFFFFFF1;
    // rom_array[24582] = 32'hFFFFFFF1;
    // rom_array[24583] = 32'hFFFFFFF1;
    // rom_array[24584] = 32'hFFFFFFF1;
    // rom_array[24585] = 32'hFFFFFFF0;
    // rom_array[24586] = 32'hFFFFFFF0;
    // rom_array[24587] = 32'hFFFFFFF0;
    // rom_array[24588] = 32'hFFFFFFF0;
    // rom_array[24589] = 32'hFFFFFFF1;
    // rom_array[24590] = 32'hFFFFFFF1;
    // rom_array[24591] = 32'hFFFFFFF1;
    // rom_array[24592] = 32'hFFFFFFF1;
    // rom_array[24593] = 32'hFFFFFFF0;
    // rom_array[24594] = 32'hFFFFFFF0;
    // rom_array[24595] = 32'hFFFFFFF0;
    // rom_array[24596] = 32'hFFFFFFF0;
    // rom_array[24597] = 32'hFFFFFFF1;
    // rom_array[24598] = 32'hFFFFFFF1;
    // rom_array[24599] = 32'hFFFFFFF1;
    // rom_array[24600] = 32'hFFFFFFF1;
    // rom_array[24601] = 32'hFFFFFFF0;
    // rom_array[24602] = 32'hFFFFFFF0;
    // rom_array[24603] = 32'hFFFFFFF0;
    // rom_array[24604] = 32'hFFFFFFF0;
    // rom_array[24605] = 32'hFFFFFFF1;
    // rom_array[24606] = 32'hFFFFFFF1;
    // rom_array[24607] = 32'hFFFFFFF1;
    // rom_array[24608] = 32'hFFFFFFF1;
    // rom_array[24609] = 32'hFFFFFFF0;
    // rom_array[24610] = 32'hFFFFFFF0;
    // rom_array[24611] = 32'hFFFFFFF0;
    // rom_array[24612] = 32'hFFFFFFF0;
    // rom_array[24613] = 32'hFFFFFFF1;
    // rom_array[24614] = 32'hFFFFFFF1;
    // rom_array[24615] = 32'hFFFFFFF1;
    // rom_array[24616] = 32'hFFFFFFF1;
    // rom_array[24617] = 32'hFFFFFFF0;
    // rom_array[24618] = 32'hFFFFFFF0;
    // rom_array[24619] = 32'hFFFFFFF0;
    // rom_array[24620] = 32'hFFFFFFF0;
    // rom_array[24621] = 32'hFFFFFFF1;
    // rom_array[24622] = 32'hFFFFFFF1;
    // rom_array[24623] = 32'hFFFFFFF1;
    // rom_array[24624] = 32'hFFFFFFF1;
    // rom_array[24625] = 32'hFFFFFFF0;
    // rom_array[24626] = 32'hFFFFFFF0;
    // rom_array[24627] = 32'hFFFFFFF0;
    // rom_array[24628] = 32'hFFFFFFF0;
    // rom_array[24629] = 32'hFFFFFFF1;
    // rom_array[24630] = 32'hFFFFFFF1;
    // rom_array[24631] = 32'hFFFFFFF1;
    // rom_array[24632] = 32'hFFFFFFF1;
    // rom_array[24633] = 32'hFFFFFFF0;
    // rom_array[24634] = 32'hFFFFFFF0;
    // rom_array[24635] = 32'hFFFFFFF0;
    // rom_array[24636] = 32'hFFFFFFF0;
    // rom_array[24637] = 32'hFFFFFFF1;
    // rom_array[24638] = 32'hFFFFFFF1;
    // rom_array[24639] = 32'hFFFFFFF1;
    // rom_array[24640] = 32'hFFFFFFF1;
    // rom_array[24641] = 32'hFFFFFFF0;
    // rom_array[24642] = 32'hFFFFFFF0;
    // rom_array[24643] = 32'hFFFFFFF0;
    // rom_array[24644] = 32'hFFFFFFF0;
    // rom_array[24645] = 32'hFFFFFFF1;
    // rom_array[24646] = 32'hFFFFFFF1;
    // rom_array[24647] = 32'hFFFFFFF1;
    // rom_array[24648] = 32'hFFFFFFF1;
    // rom_array[24649] = 32'hFFFFFFF1;
    // rom_array[24650] = 32'hFFFFFFF1;
    // rom_array[24651] = 32'hFFFFFFF1;
    // rom_array[24652] = 32'hFFFFFFF1;
    // rom_array[24653] = 32'hFFFFFFF1;
    // rom_array[24654] = 32'hFFFFFFF1;
    // rom_array[24655] = 32'hFFFFFFF1;
    // rom_array[24656] = 32'hFFFFFFF1;
    // rom_array[24657] = 32'hFFFFFFF1;
    // rom_array[24658] = 32'hFFFFFFF1;
    // rom_array[24659] = 32'hFFFFFFF1;
    // rom_array[24660] = 32'hFFFFFFF1;
    // rom_array[24661] = 32'hFFFFFFF1;
    // rom_array[24662] = 32'hFFFFFFF1;
    // rom_array[24663] = 32'hFFFFFFF1;
    // rom_array[24664] = 32'hFFFFFFF1;
    // rom_array[24665] = 32'hFFFFFFF1;
    // rom_array[24666] = 32'hFFFFFFF1;
    // rom_array[24667] = 32'hFFFFFFF1;
    // rom_array[24668] = 32'hFFFFFFF1;
    // rom_array[24669] = 32'hFFFFFFF1;
    // rom_array[24670] = 32'hFFFFFFF1;
    // rom_array[24671] = 32'hFFFFFFF1;
    // rom_array[24672] = 32'hFFFFFFF1;
    // rom_array[24673] = 32'hFFFFFFF1;
    // rom_array[24674] = 32'hFFFFFFF1;
    // rom_array[24675] = 32'hFFFFFFF1;
    // rom_array[24676] = 32'hFFFFFFF1;
    // rom_array[24677] = 32'hFFFFFFF1;
    // rom_array[24678] = 32'hFFFFFFF1;
    // rom_array[24679] = 32'hFFFFFFF1;
    // rom_array[24680] = 32'hFFFFFFF1;
    // rom_array[24681] = 32'hFFFFFFF1;
    // rom_array[24682] = 32'hFFFFFFF1;
    // rom_array[24683] = 32'hFFFFFFF1;
    // rom_array[24684] = 32'hFFFFFFF1;
    // rom_array[24685] = 32'hFFFFFFF1;
    // rom_array[24686] = 32'hFFFFFFF1;
    // rom_array[24687] = 32'hFFFFFFF1;
    // rom_array[24688] = 32'hFFFFFFF1;
    // rom_array[24689] = 32'hFFFFFFF1;
    // rom_array[24690] = 32'hFFFFFFF1;
    // rom_array[24691] = 32'hFFFFFFF1;
    // rom_array[24692] = 32'hFFFFFFF1;
    // rom_array[24693] = 32'hFFFFFFF1;
    // rom_array[24694] = 32'hFFFFFFF1;
    // rom_array[24695] = 32'hFFFFFFF1;
    // rom_array[24696] = 32'hFFFFFFF1;
    // rom_array[24697] = 32'hFFFFFFF1;
    // rom_array[24698] = 32'hFFFFFFF1;
    // rom_array[24699] = 32'hFFFFFFF1;
    // rom_array[24700] = 32'hFFFFFFF1;
    // rom_array[24701] = 32'hFFFFFFF0;
    // rom_array[24702] = 32'hFFFFFFF0;
    // rom_array[24703] = 32'hFFFFFFF0;
    // rom_array[24704] = 32'hFFFFFFF0;
    // rom_array[24705] = 32'hFFFFFFF1;
    // rom_array[24706] = 32'hFFFFFFF1;
    // rom_array[24707] = 32'hFFFFFFF1;
    // rom_array[24708] = 32'hFFFFFFF1;
    // rom_array[24709] = 32'hFFFFFFF0;
    // rom_array[24710] = 32'hFFFFFFF0;
    // rom_array[24711] = 32'hFFFFFFF0;
    // rom_array[24712] = 32'hFFFFFFF0;
    // rom_array[24713] = 32'hFFFFFFF1;
    // rom_array[24714] = 32'hFFFFFFF1;
    // rom_array[24715] = 32'hFFFFFFF1;
    // rom_array[24716] = 32'hFFFFFFF1;
    // rom_array[24717] = 32'hFFFFFFF0;
    // rom_array[24718] = 32'hFFFFFFF0;
    // rom_array[24719] = 32'hFFFFFFF0;
    // rom_array[24720] = 32'hFFFFFFF0;
    // rom_array[24721] = 32'hFFFFFFF1;
    // rom_array[24722] = 32'hFFFFFFF1;
    // rom_array[24723] = 32'hFFFFFFF1;
    // rom_array[24724] = 32'hFFFFFFF1;
    // rom_array[24725] = 32'hFFFFFFF0;
    // rom_array[24726] = 32'hFFFFFFF0;
    // rom_array[24727] = 32'hFFFFFFF0;
    // rom_array[24728] = 32'hFFFFFFF0;
    // rom_array[24729] = 32'hFFFFFFF1;
    // rom_array[24730] = 32'hFFFFFFF1;
    // rom_array[24731] = 32'hFFFFFFF1;
    // rom_array[24732] = 32'hFFFFFFF1;
    // rom_array[24733] = 32'hFFFFFFF0;
    // rom_array[24734] = 32'hFFFFFFF0;
    // rom_array[24735] = 32'hFFFFFFF0;
    // rom_array[24736] = 32'hFFFFFFF0;
    // rom_array[24737] = 32'hFFFFFFF1;
    // rom_array[24738] = 32'hFFFFFFF1;
    // rom_array[24739] = 32'hFFFFFFF1;
    // rom_array[24740] = 32'hFFFFFFF1;
    // rom_array[24741] = 32'hFFFFFFF0;
    // rom_array[24742] = 32'hFFFFFFF0;
    // rom_array[24743] = 32'hFFFFFFF0;
    // rom_array[24744] = 32'hFFFFFFF0;
    // rom_array[24745] = 32'hFFFFFFF1;
    // rom_array[24746] = 32'hFFFFFFF1;
    // rom_array[24747] = 32'hFFFFFFF1;
    // rom_array[24748] = 32'hFFFFFFF1;
    // rom_array[24749] = 32'hFFFFFFF0;
    // rom_array[24750] = 32'hFFFFFFF0;
    // rom_array[24751] = 32'hFFFFFFF0;
    // rom_array[24752] = 32'hFFFFFFF0;
    // rom_array[24753] = 32'hFFFFFFF1;
    // rom_array[24754] = 32'hFFFFFFF1;
    // rom_array[24755] = 32'hFFFFFFF1;
    // rom_array[24756] = 32'hFFFFFFF1;
    // rom_array[24757] = 32'hFFFFFFF0;
    // rom_array[24758] = 32'hFFFFFFF0;
    // rom_array[24759] = 32'hFFFFFFF0;
    // rom_array[24760] = 32'hFFFFFFF0;
    // rom_array[24761] = 32'hFFFFFFF1;
    // rom_array[24762] = 32'hFFFFFFF1;
    // rom_array[24763] = 32'hFFFFFFF1;
    // rom_array[24764] = 32'hFFFFFFF1;
    // rom_array[24765] = 32'hFFFFFFF0;
    // rom_array[24766] = 32'hFFFFFFF0;
    // rom_array[24767] = 32'hFFFFFFF1;
    // rom_array[24768] = 32'hFFFFFFF1;
    // rom_array[24769] = 32'hFFFFFFF1;
    // rom_array[24770] = 32'hFFFFFFF1;
    // rom_array[24771] = 32'hFFFFFFF1;
    // rom_array[24772] = 32'hFFFFFFF1;
    // rom_array[24773] = 32'hFFFFFFF0;
    // rom_array[24774] = 32'hFFFFFFF0;
    // rom_array[24775] = 32'hFFFFFFF1;
    // rom_array[24776] = 32'hFFFFFFF1;
    // rom_array[24777] = 32'hFFFFFFF1;
    // rom_array[24778] = 32'hFFFFFFF1;
    // rom_array[24779] = 32'hFFFFFFF1;
    // rom_array[24780] = 32'hFFFFFFF1;
    // rom_array[24781] = 32'hFFFFFFF1;
    // rom_array[24782] = 32'hFFFFFFF1;
    // rom_array[24783] = 32'hFFFFFFF1;
    // rom_array[24784] = 32'hFFFFFFF1;
    // rom_array[24785] = 32'hFFFFFFF1;
    // rom_array[24786] = 32'hFFFFFFF1;
    // rom_array[24787] = 32'hFFFFFFF1;
    // rom_array[24788] = 32'hFFFFFFF1;
    // rom_array[24789] = 32'hFFFFFFF1;
    // rom_array[24790] = 32'hFFFFFFF1;
    // rom_array[24791] = 32'hFFFFFFF1;
    // rom_array[24792] = 32'hFFFFFFF1;
    // rom_array[24793] = 32'hFFFFFFF0;
    // rom_array[24794] = 32'hFFFFFFF0;
    // rom_array[24795] = 32'hFFFFFFF1;
    // rom_array[24796] = 32'hFFFFFFF1;
    // rom_array[24797] = 32'hFFFFFFF0;
    // rom_array[24798] = 32'hFFFFFFF0;
    // rom_array[24799] = 32'hFFFFFFF1;
    // rom_array[24800] = 32'hFFFFFFF1;
    // rom_array[24801] = 32'hFFFFFFF0;
    // rom_array[24802] = 32'hFFFFFFF0;
    // rom_array[24803] = 32'hFFFFFFF1;
    // rom_array[24804] = 32'hFFFFFFF1;
    // rom_array[24805] = 32'hFFFFFFF0;
    // rom_array[24806] = 32'hFFFFFFF0;
    // rom_array[24807] = 32'hFFFFFFF1;
    // rom_array[24808] = 32'hFFFFFFF1;
    // rom_array[24809] = 32'hFFFFFFF0;
    // rom_array[24810] = 32'hFFFFFFF0;
    // rom_array[24811] = 32'hFFFFFFF0;
    // rom_array[24812] = 32'hFFFFFFF0;
    // rom_array[24813] = 32'hFFFFFFF1;
    // rom_array[24814] = 32'hFFFFFFF1;
    // rom_array[24815] = 32'hFFFFFFF1;
    // rom_array[24816] = 32'hFFFFFFF1;
    // rom_array[24817] = 32'hFFFFFFF0;
    // rom_array[24818] = 32'hFFFFFFF0;
    // rom_array[24819] = 32'hFFFFFFF0;
    // rom_array[24820] = 32'hFFFFFFF0;
    // rom_array[24821] = 32'hFFFFFFF1;
    // rom_array[24822] = 32'hFFFFFFF1;
    // rom_array[24823] = 32'hFFFFFFF1;
    // rom_array[24824] = 32'hFFFFFFF1;
    // rom_array[24825] = 32'hFFFFFFF0;
    // rom_array[24826] = 32'hFFFFFFF0;
    // rom_array[24827] = 32'hFFFFFFF0;
    // rom_array[24828] = 32'hFFFFFFF0;
    // rom_array[24829] = 32'hFFFFFFF1;
    // rom_array[24830] = 32'hFFFFFFF1;
    // rom_array[24831] = 32'hFFFFFFF1;
    // rom_array[24832] = 32'hFFFFFFF1;
    // rom_array[24833] = 32'hFFFFFFF0;
    // rom_array[24834] = 32'hFFFFFFF0;
    // rom_array[24835] = 32'hFFFFFFF0;
    // rom_array[24836] = 32'hFFFFFFF0;
    // rom_array[24837] = 32'hFFFFFFF1;
    // rom_array[24838] = 32'hFFFFFFF1;
    // rom_array[24839] = 32'hFFFFFFF1;
    // rom_array[24840] = 32'hFFFFFFF1;
    // rom_array[24841] = 32'hFFFFFFF0;
    // rom_array[24842] = 32'hFFFFFFF0;
    // rom_array[24843] = 32'hFFFFFFF0;
    // rom_array[24844] = 32'hFFFFFFF0;
    // rom_array[24845] = 32'hFFFFFFF1;
    // rom_array[24846] = 32'hFFFFFFF1;
    // rom_array[24847] = 32'hFFFFFFF1;
    // rom_array[24848] = 32'hFFFFFFF1;
    // rom_array[24849] = 32'hFFFFFFF0;
    // rom_array[24850] = 32'hFFFFFFF0;
    // rom_array[24851] = 32'hFFFFFFF0;
    // rom_array[24852] = 32'hFFFFFFF0;
    // rom_array[24853] = 32'hFFFFFFF1;
    // rom_array[24854] = 32'hFFFFFFF1;
    // rom_array[24855] = 32'hFFFFFFF1;
    // rom_array[24856] = 32'hFFFFFFF1;
    // rom_array[24857] = 32'hFFFFFFF1;
    // rom_array[24858] = 32'hFFFFFFF1;
    // rom_array[24859] = 32'hFFFFFFF1;
    // rom_array[24860] = 32'hFFFFFFF1;
    // rom_array[24861] = 32'hFFFFFFF1;
    // rom_array[24862] = 32'hFFFFFFF1;
    // rom_array[24863] = 32'hFFFFFFF1;
    // rom_array[24864] = 32'hFFFFFFF1;
    // rom_array[24865] = 32'hFFFFFFF1;
    // rom_array[24866] = 32'hFFFFFFF1;
    // rom_array[24867] = 32'hFFFFFFF1;
    // rom_array[24868] = 32'hFFFFFFF1;
    // rom_array[24869] = 32'hFFFFFFF1;
    // rom_array[24870] = 32'hFFFFFFF1;
    // rom_array[24871] = 32'hFFFFFFF1;
    // rom_array[24872] = 32'hFFFFFFF1;
    // rom_array[24873] = 32'hFFFFFFF1;
    // rom_array[24874] = 32'hFFFFFFF1;
    // rom_array[24875] = 32'hFFFFFFF1;
    // rom_array[24876] = 32'hFFFFFFF1;
    // rom_array[24877] = 32'hFFFFFFF1;
    // rom_array[24878] = 32'hFFFFFFF1;
    // rom_array[24879] = 32'hFFFFFFF1;
    // rom_array[24880] = 32'hFFFFFFF1;
    // rom_array[24881] = 32'hFFFFFFF1;
    // rom_array[24882] = 32'hFFFFFFF1;
    // rom_array[24883] = 32'hFFFFFFF1;
    // rom_array[24884] = 32'hFFFFFFF1;
    // rom_array[24885] = 32'hFFFFFFF1;
    // rom_array[24886] = 32'hFFFFFFF1;
    // rom_array[24887] = 32'hFFFFFFF1;
    // rom_array[24888] = 32'hFFFFFFF1;
    // rom_array[24889] = 32'hFFFFFFF1;
    // rom_array[24890] = 32'hFFFFFFF1;
    // rom_array[24891] = 32'hFFFFFFF1;
    // rom_array[24892] = 32'hFFFFFFF1;
    // rom_array[24893] = 32'hFFFFFFF1;
    // rom_array[24894] = 32'hFFFFFFF1;
    // rom_array[24895] = 32'hFFFFFFF1;
    // rom_array[24896] = 32'hFFFFFFF1;
    // rom_array[24897] = 32'hFFFFFFF1;
    // rom_array[24898] = 32'hFFFFFFF1;
    // rom_array[24899] = 32'hFFFFFFF1;
    // rom_array[24900] = 32'hFFFFFFF1;
    // rom_array[24901] = 32'hFFFFFFF1;
    // rom_array[24902] = 32'hFFFFFFF1;
    // rom_array[24903] = 32'hFFFFFFF1;
    // rom_array[24904] = 32'hFFFFFFF1;
    // rom_array[24905] = 32'hFFFFFFF1;
    // rom_array[24906] = 32'hFFFFFFF1;
    // rom_array[24907] = 32'hFFFFFFF1;
    // rom_array[24908] = 32'hFFFFFFF1;
    // rom_array[24909] = 32'hFFFFFFF1;
    // rom_array[24910] = 32'hFFFFFFF1;
    // rom_array[24911] = 32'hFFFFFFF1;
    // rom_array[24912] = 32'hFFFFFFF1;
    // rom_array[24913] = 32'hFFFFFFF1;
    // rom_array[24914] = 32'hFFFFFFF1;
    // rom_array[24915] = 32'hFFFFFFF1;
    // rom_array[24916] = 32'hFFFFFFF1;
    // rom_array[24917] = 32'hFFFFFFF1;
    // rom_array[24918] = 32'hFFFFFFF1;
    // rom_array[24919] = 32'hFFFFFFF1;
    // rom_array[24920] = 32'hFFFFFFF1;
    // rom_array[24921] = 32'hFFFFFFF1;
    // rom_array[24922] = 32'hFFFFFFF1;
    // rom_array[24923] = 32'hFFFFFFF1;
    // rom_array[24924] = 32'hFFFFFFF1;
    // rom_array[24925] = 32'hFFFFFFF1;
    // rom_array[24926] = 32'hFFFFFFF1;
    // rom_array[24927] = 32'hFFFFFFF1;
    // rom_array[24928] = 32'hFFFFFFF1;
    // rom_array[24929] = 32'hFFFFFFF1;
    // rom_array[24930] = 32'hFFFFFFF1;
    // rom_array[24931] = 32'hFFFFFFF1;
    // rom_array[24932] = 32'hFFFFFFF1;
    // rom_array[24933] = 32'hFFFFFFF1;
    // rom_array[24934] = 32'hFFFFFFF1;
    // rom_array[24935] = 32'hFFFFFFF1;
    // rom_array[24936] = 32'hFFFFFFF1;
    // rom_array[24937] = 32'hFFFFFFF1;
    // rom_array[24938] = 32'hFFFFFFF1;
    // rom_array[24939] = 32'hFFFFFFF1;
    // rom_array[24940] = 32'hFFFFFFF1;
    // rom_array[24941] = 32'hFFFFFFF1;
    // rom_array[24942] = 32'hFFFFFFF1;
    // rom_array[24943] = 32'hFFFFFFF1;
    // rom_array[24944] = 32'hFFFFFFF1;
    // rom_array[24945] = 32'hFFFFFFF1;
    // rom_array[24946] = 32'hFFFFFFF1;
    // rom_array[24947] = 32'hFFFFFFF1;
    // rom_array[24948] = 32'hFFFFFFF1;
    // rom_array[24949] = 32'hFFFFFFF1;
    // rom_array[24950] = 32'hFFFFFFF1;
    // rom_array[24951] = 32'hFFFFFFF1;
    // rom_array[24952] = 32'hFFFFFFF1;
    // rom_array[24953] = 32'hFFFFFFF1;
    // rom_array[24954] = 32'hFFFFFFF1;
    // rom_array[24955] = 32'hFFFFFFF1;
    // rom_array[24956] = 32'hFFFFFFF1;
    // rom_array[24957] = 32'hFFFFFFF1;
    // rom_array[24958] = 32'hFFFFFFF1;
    // rom_array[24959] = 32'hFFFFFFF1;
    // rom_array[24960] = 32'hFFFFFFF1;
    // rom_array[24961] = 32'hFFFFFFF1;
    // rom_array[24962] = 32'hFFFFFFF1;
    // rom_array[24963] = 32'hFFFFFFF1;
    // rom_array[24964] = 32'hFFFFFFF1;
    // rom_array[24965] = 32'hFFFFFFF1;
    // rom_array[24966] = 32'hFFFFFFF1;
    // rom_array[24967] = 32'hFFFFFFF1;
    // rom_array[24968] = 32'hFFFFFFF1;
    // rom_array[24969] = 32'hFFFFFFF1;
    // rom_array[24970] = 32'hFFFFFFF1;
    // rom_array[24971] = 32'hFFFFFFF1;
    // rom_array[24972] = 32'hFFFFFFF1;
    // rom_array[24973] = 32'hFFFFFFF1;
    // rom_array[24974] = 32'hFFFFFFF1;
    // rom_array[24975] = 32'hFFFFFFF1;
    // rom_array[24976] = 32'hFFFFFFF1;
    // rom_array[24977] = 32'hFFFFFFF1;
    // rom_array[24978] = 32'hFFFFFFF1;
    // rom_array[24979] = 32'hFFFFFFF1;
    // rom_array[24980] = 32'hFFFFFFF1;
    // rom_array[24981] = 32'hFFFFFFF1;
    // rom_array[24982] = 32'hFFFFFFF1;
    // rom_array[24983] = 32'hFFFFFFF1;
    // rom_array[24984] = 32'hFFFFFFF1;
    // rom_array[24985] = 32'hFFFFFFF1;
    // rom_array[24986] = 32'hFFFFFFF1;
    // rom_array[24987] = 32'hFFFFFFF1;
    // rom_array[24988] = 32'hFFFFFFF1;
    // rom_array[24989] = 32'hFFFFFFF1;
    // rom_array[24990] = 32'hFFFFFFF1;
    // rom_array[24991] = 32'hFFFFFFF1;
    // rom_array[24992] = 32'hFFFFFFF1;
    // rom_array[24993] = 32'hFFFFFFF1;
    // rom_array[24994] = 32'hFFFFFFF1;
    // rom_array[24995] = 32'hFFFFFFF1;
    // rom_array[24996] = 32'hFFFFFFF1;
    // rom_array[24997] = 32'hFFFFFFF1;
    // rom_array[24998] = 32'hFFFFFFF1;
    // rom_array[24999] = 32'hFFFFFFF1;
    // rom_array[25000] = 32'hFFFFFFF1;
    // rom_array[25001] = 32'hFFFFFFF1;
    // rom_array[25002] = 32'hFFFFFFF1;
    // rom_array[25003] = 32'hFFFFFFF1;
    // rom_array[25004] = 32'hFFFFFFF1;
    // rom_array[25005] = 32'hFFFFFFF1;
    // rom_array[25006] = 32'hFFFFFFF1;
    // rom_array[25007] = 32'hFFFFFFF1;
    // rom_array[25008] = 32'hFFFFFFF1;
    // rom_array[25009] = 32'hFFFFFFF1;
    // rom_array[25010] = 32'hFFFFFFF1;
    // rom_array[25011] = 32'hFFFFFFF1;
    // rom_array[25012] = 32'hFFFFFFF1;
    // rom_array[25013] = 32'hFFFFFFF1;
    // rom_array[25014] = 32'hFFFFFFF1;
    // rom_array[25015] = 32'hFFFFFFF1;
    // rom_array[25016] = 32'hFFFFFFF1;
    // rom_array[25017] = 32'hFFFFFFF1;
    // rom_array[25018] = 32'hFFFFFFF1;
    // rom_array[25019] = 32'hFFFFFFF1;
    // rom_array[25020] = 32'hFFFFFFF1;
    // rom_array[25021] = 32'hFFFFFFF1;
    // rom_array[25022] = 32'hFFFFFFF1;
    // rom_array[25023] = 32'hFFFFFFF1;
    // rom_array[25024] = 32'hFFFFFFF1;
    // rom_array[25025] = 32'hFFFFFFF1;
    // rom_array[25026] = 32'hFFFFFFF1;
    // rom_array[25027] = 32'hFFFFFFF1;
    // rom_array[25028] = 32'hFFFFFFF1;
    // rom_array[25029] = 32'hFFFFFFF1;
    // rom_array[25030] = 32'hFFFFFFF1;
    // rom_array[25031] = 32'hFFFFFFF1;
    // rom_array[25032] = 32'hFFFFFFF1;
    // rom_array[25033] = 32'hFFFFFFF0;
    // rom_array[25034] = 32'hFFFFFFF0;
    // rom_array[25035] = 32'hFFFFFFF1;
    // rom_array[25036] = 32'hFFFFFFF1;
    // rom_array[25037] = 32'hFFFFFFF0;
    // rom_array[25038] = 32'hFFFFFFF0;
    // rom_array[25039] = 32'hFFFFFFF1;
    // rom_array[25040] = 32'hFFFFFFF1;
    // rom_array[25041] = 32'hFFFFFFF0;
    // rom_array[25042] = 32'hFFFFFFF0;
    // rom_array[25043] = 32'hFFFFFFF1;
    // rom_array[25044] = 32'hFFFFFFF1;
    // rom_array[25045] = 32'hFFFFFFF0;
    // rom_array[25046] = 32'hFFFFFFF0;
    // rom_array[25047] = 32'hFFFFFFF1;
    // rom_array[25048] = 32'hFFFFFFF1;
    // rom_array[25049] = 32'hFFFFFFF0;
    // rom_array[25050] = 32'hFFFFFFF0;
    // rom_array[25051] = 32'hFFFFFFF1;
    // rom_array[25052] = 32'hFFFFFFF1;
    // rom_array[25053] = 32'hFFFFFFF0;
    // rom_array[25054] = 32'hFFFFFFF0;
    // rom_array[25055] = 32'hFFFFFFF1;
    // rom_array[25056] = 32'hFFFFFFF1;
    // rom_array[25057] = 32'hFFFFFFF0;
    // rom_array[25058] = 32'hFFFFFFF0;
    // rom_array[25059] = 32'hFFFFFFF1;
    // rom_array[25060] = 32'hFFFFFFF1;
    // rom_array[25061] = 32'hFFFFFFF0;
    // rom_array[25062] = 32'hFFFFFFF0;
    // rom_array[25063] = 32'hFFFFFFF1;
    // rom_array[25064] = 32'hFFFFFFF1;
    // rom_array[25065] = 32'hFFFFFFF0;
    // rom_array[25066] = 32'hFFFFFFF0;
    // rom_array[25067] = 32'hFFFFFFF1;
    // rom_array[25068] = 32'hFFFFFFF1;
    // rom_array[25069] = 32'hFFFFFFF0;
    // rom_array[25070] = 32'hFFFFFFF0;
    // rom_array[25071] = 32'hFFFFFFF1;
    // rom_array[25072] = 32'hFFFFFFF1;
    // rom_array[25073] = 32'hFFFFFFF0;
    // rom_array[25074] = 32'hFFFFFFF0;
    // rom_array[25075] = 32'hFFFFFFF1;
    // rom_array[25076] = 32'hFFFFFFF1;
    // rom_array[25077] = 32'hFFFFFFF0;
    // rom_array[25078] = 32'hFFFFFFF0;
    // rom_array[25079] = 32'hFFFFFFF1;
    // rom_array[25080] = 32'hFFFFFFF1;
    // rom_array[25081] = 32'hFFFFFFF0;
    // rom_array[25082] = 32'hFFFFFFF0;
    // rom_array[25083] = 32'hFFFFFFF1;
    // rom_array[25084] = 32'hFFFFFFF1;
    // rom_array[25085] = 32'hFFFFFFF0;
    // rom_array[25086] = 32'hFFFFFFF0;
    // rom_array[25087] = 32'hFFFFFFF1;
    // rom_array[25088] = 32'hFFFFFFF1;
    // rom_array[25089] = 32'hFFFFFFF0;
    // rom_array[25090] = 32'hFFFFFFF0;
    // rom_array[25091] = 32'hFFFFFFF1;
    // rom_array[25092] = 32'hFFFFFFF1;
    // rom_array[25093] = 32'hFFFFFFF0;
    // rom_array[25094] = 32'hFFFFFFF0;
    // rom_array[25095] = 32'hFFFFFFF1;
    // rom_array[25096] = 32'hFFFFFFF1;
    // rom_array[25097] = 32'hFFFFFFF1;
    // rom_array[25098] = 32'hFFFFFFF1;
    // rom_array[25099] = 32'hFFFFFFF1;
    // rom_array[25100] = 32'hFFFFFFF1;
    // rom_array[25101] = 32'hFFFFFFF1;
    // rom_array[25102] = 32'hFFFFFFF1;
    // rom_array[25103] = 32'hFFFFFFF1;
    // rom_array[25104] = 32'hFFFFFFF1;
    // rom_array[25105] = 32'hFFFFFFF1;
    // rom_array[25106] = 32'hFFFFFFF1;
    // rom_array[25107] = 32'hFFFFFFF1;
    // rom_array[25108] = 32'hFFFFFFF1;
    // rom_array[25109] = 32'hFFFFFFF1;
    // rom_array[25110] = 32'hFFFFFFF1;
    // rom_array[25111] = 32'hFFFFFFF1;
    // rom_array[25112] = 32'hFFFFFFF1;
    // rom_array[25113] = 32'hFFFFFFF1;
    // rom_array[25114] = 32'hFFFFFFF1;
    // rom_array[25115] = 32'hFFFFFFF1;
    // rom_array[25116] = 32'hFFFFFFF1;
    // rom_array[25117] = 32'hFFFFFFF1;
    // rom_array[25118] = 32'hFFFFFFF1;
    // rom_array[25119] = 32'hFFFFFFF1;
    // rom_array[25120] = 32'hFFFFFFF1;
    // rom_array[25121] = 32'hFFFFFFF1;
    // rom_array[25122] = 32'hFFFFFFF1;
    // rom_array[25123] = 32'hFFFFFFF1;
    // rom_array[25124] = 32'hFFFFFFF1;
    // rom_array[25125] = 32'hFFFFFFF1;
    // rom_array[25126] = 32'hFFFFFFF1;
    // rom_array[25127] = 32'hFFFFFFF1;
    // rom_array[25128] = 32'hFFFFFFF1;
    // rom_array[25129] = 32'hFFFFFFF1;
    // rom_array[25130] = 32'hFFFFFFF1;
    // rom_array[25131] = 32'hFFFFFFF1;
    // rom_array[25132] = 32'hFFFFFFF1;
    // rom_array[25133] = 32'hFFFFFFF1;
    // rom_array[25134] = 32'hFFFFFFF1;
    // rom_array[25135] = 32'hFFFFFFF1;
    // rom_array[25136] = 32'hFFFFFFF1;
    // rom_array[25137] = 32'hFFFFFFF1;
    // rom_array[25138] = 32'hFFFFFFF1;
    // rom_array[25139] = 32'hFFFFFFF1;
    // rom_array[25140] = 32'hFFFFFFF1;
    // rom_array[25141] = 32'hFFFFFFF1;
    // rom_array[25142] = 32'hFFFFFFF1;
    // rom_array[25143] = 32'hFFFFFFF1;
    // rom_array[25144] = 32'hFFFFFFF1;
    // rom_array[25145] = 32'hFFFFFFF1;
    // rom_array[25146] = 32'hFFFFFFF1;
    // rom_array[25147] = 32'hFFFFFFF1;
    // rom_array[25148] = 32'hFFFFFFF1;
    // rom_array[25149] = 32'hFFFFFFF1;
    // rom_array[25150] = 32'hFFFFFFF1;
    // rom_array[25151] = 32'hFFFFFFF1;
    // rom_array[25152] = 32'hFFFFFFF1;
    // rom_array[25153] = 32'hFFFFFFF1;
    // rom_array[25154] = 32'hFFFFFFF1;
    // rom_array[25155] = 32'hFFFFFFF1;
    // rom_array[25156] = 32'hFFFFFFF1;
    // rom_array[25157] = 32'hFFFFFFF1;
    // rom_array[25158] = 32'hFFFFFFF1;
    // rom_array[25159] = 32'hFFFFFFF1;
    // rom_array[25160] = 32'hFFFFFFF1;
    // rom_array[25161] = 32'hFFFFFFF0;
    // rom_array[25162] = 32'hFFFFFFF0;
    // rom_array[25163] = 32'hFFFFFFF1;
    // rom_array[25164] = 32'hFFFFFFF1;
    // rom_array[25165] = 32'hFFFFFFF0;
    // rom_array[25166] = 32'hFFFFFFF0;
    // rom_array[25167] = 32'hFFFFFFF1;
    // rom_array[25168] = 32'hFFFFFFF1;
    // rom_array[25169] = 32'hFFFFFFF0;
    // rom_array[25170] = 32'hFFFFFFF0;
    // rom_array[25171] = 32'hFFFFFFF1;
    // rom_array[25172] = 32'hFFFFFFF1;
    // rom_array[25173] = 32'hFFFFFFF0;
    // rom_array[25174] = 32'hFFFFFFF0;
    // rom_array[25175] = 32'hFFFFFFF1;
    // rom_array[25176] = 32'hFFFFFFF1;
    // rom_array[25177] = 32'hFFFFFFF0;
    // rom_array[25178] = 32'hFFFFFFF0;
    // rom_array[25179] = 32'hFFFFFFF1;
    // rom_array[25180] = 32'hFFFFFFF1;
    // rom_array[25181] = 32'hFFFFFFF0;
    // rom_array[25182] = 32'hFFFFFFF0;
    // rom_array[25183] = 32'hFFFFFFF1;
    // rom_array[25184] = 32'hFFFFFFF1;
    // rom_array[25185] = 32'hFFFFFFF0;
    // rom_array[25186] = 32'hFFFFFFF0;
    // rom_array[25187] = 32'hFFFFFFF1;
    // rom_array[25188] = 32'hFFFFFFF1;
    // rom_array[25189] = 32'hFFFFFFF0;
    // rom_array[25190] = 32'hFFFFFFF0;
    // rom_array[25191] = 32'hFFFFFFF1;
    // rom_array[25192] = 32'hFFFFFFF1;
    // rom_array[25193] = 32'hFFFFFFF0;
    // rom_array[25194] = 32'hFFFFFFF0;
    // rom_array[25195] = 32'hFFFFFFF1;
    // rom_array[25196] = 32'hFFFFFFF1;
    // rom_array[25197] = 32'hFFFFFFF0;
    // rom_array[25198] = 32'hFFFFFFF0;
    // rom_array[25199] = 32'hFFFFFFF1;
    // rom_array[25200] = 32'hFFFFFFF1;
    // rom_array[25201] = 32'hFFFFFFF0;
    // rom_array[25202] = 32'hFFFFFFF0;
    // rom_array[25203] = 32'hFFFFFFF1;
    // rom_array[25204] = 32'hFFFFFFF1;
    // rom_array[25205] = 32'hFFFFFFF0;
    // rom_array[25206] = 32'hFFFFFFF0;
    // rom_array[25207] = 32'hFFFFFFF1;
    // rom_array[25208] = 32'hFFFFFFF1;
    // rom_array[25209] = 32'hFFFFFFF0;
    // rom_array[25210] = 32'hFFFFFFF0;
    // rom_array[25211] = 32'hFFFFFFF1;
    // rom_array[25212] = 32'hFFFFFFF1;
    // rom_array[25213] = 32'hFFFFFFF0;
    // rom_array[25214] = 32'hFFFFFFF0;
    // rom_array[25215] = 32'hFFFFFFF1;
    // rom_array[25216] = 32'hFFFFFFF1;
    // rom_array[25217] = 32'hFFFFFFF0;
    // rom_array[25218] = 32'hFFFFFFF0;
    // rom_array[25219] = 32'hFFFFFFF1;
    // rom_array[25220] = 32'hFFFFFFF1;
    // rom_array[25221] = 32'hFFFFFFF0;
    // rom_array[25222] = 32'hFFFFFFF0;
    // rom_array[25223] = 32'hFFFFFFF1;
    // rom_array[25224] = 32'hFFFFFFF1;
    // rom_array[25225] = 32'hFFFFFFF1;
    // rom_array[25226] = 32'hFFFFFFF1;
    // rom_array[25227] = 32'hFFFFFFF1;
    // rom_array[25228] = 32'hFFFFFFF1;
    // rom_array[25229] = 32'hFFFFFFF1;
    // rom_array[25230] = 32'hFFFFFFF1;
    // rom_array[25231] = 32'hFFFFFFF1;
    // rom_array[25232] = 32'hFFFFFFF1;
    // rom_array[25233] = 32'hFFFFFFF1;
    // rom_array[25234] = 32'hFFFFFFF1;
    // rom_array[25235] = 32'hFFFFFFF1;
    // rom_array[25236] = 32'hFFFFFFF1;
    // rom_array[25237] = 32'hFFFFFFF1;
    // rom_array[25238] = 32'hFFFFFFF1;
    // rom_array[25239] = 32'hFFFFFFF1;
    // rom_array[25240] = 32'hFFFFFFF1;
    // rom_array[25241] = 32'hFFFFFFF1;
    // rom_array[25242] = 32'hFFFFFFF1;
    // rom_array[25243] = 32'hFFFFFFF1;
    // rom_array[25244] = 32'hFFFFFFF1;
    // rom_array[25245] = 32'hFFFFFFF1;
    // rom_array[25246] = 32'hFFFFFFF1;
    // rom_array[25247] = 32'hFFFFFFF1;
    // rom_array[25248] = 32'hFFFFFFF1;
    // rom_array[25249] = 32'hFFFFFFF1;
    // rom_array[25250] = 32'hFFFFFFF1;
    // rom_array[25251] = 32'hFFFFFFF1;
    // rom_array[25252] = 32'hFFFFFFF1;
    // rom_array[25253] = 32'hFFFFFFF1;
    // rom_array[25254] = 32'hFFFFFFF1;
    // rom_array[25255] = 32'hFFFFFFF1;
    // rom_array[25256] = 32'hFFFFFFF1;
    // rom_array[25257] = 32'hFFFFFFF1;
    // rom_array[25258] = 32'hFFFFFFF1;
    // rom_array[25259] = 32'hFFFFFFF1;
    // rom_array[25260] = 32'hFFFFFFF1;
    // rom_array[25261] = 32'hFFFFFFF1;
    // rom_array[25262] = 32'hFFFFFFF1;
    // rom_array[25263] = 32'hFFFFFFF1;
    // rom_array[25264] = 32'hFFFFFFF1;
    // rom_array[25265] = 32'hFFFFFFF1;
    // rom_array[25266] = 32'hFFFFFFF1;
    // rom_array[25267] = 32'hFFFFFFF1;
    // rom_array[25268] = 32'hFFFFFFF1;
    // rom_array[25269] = 32'hFFFFFFF1;
    // rom_array[25270] = 32'hFFFFFFF1;
    // rom_array[25271] = 32'hFFFFFFF1;
    // rom_array[25272] = 32'hFFFFFFF1;
    // rom_array[25273] = 32'hFFFFFFF1;
    // rom_array[25274] = 32'hFFFFFFF1;
    // rom_array[25275] = 32'hFFFFFFF1;
    // rom_array[25276] = 32'hFFFFFFF1;
    // rom_array[25277] = 32'hFFFFFFF1;
    // rom_array[25278] = 32'hFFFFFFF1;
    // rom_array[25279] = 32'hFFFFFFF1;
    // rom_array[25280] = 32'hFFFFFFF1;
    // rom_array[25281] = 32'hFFFFFFF1;
    // rom_array[25282] = 32'hFFFFFFF1;
    // rom_array[25283] = 32'hFFFFFFF1;
    // rom_array[25284] = 32'hFFFFFFF1;
    // rom_array[25285] = 32'hFFFFFFF1;
    // rom_array[25286] = 32'hFFFFFFF1;
    // rom_array[25287] = 32'hFFFFFFF1;
    // rom_array[25288] = 32'hFFFFFFF1;
    // rom_array[25289] = 32'hFFFFFFF1;
    // rom_array[25290] = 32'hFFFFFFF1;
    // rom_array[25291] = 32'hFFFFFFF1;
    // rom_array[25292] = 32'hFFFFFFF1;
    // rom_array[25293] = 32'hFFFFFFF1;
    // rom_array[25294] = 32'hFFFFFFF1;
    // rom_array[25295] = 32'hFFFFFFF1;
    // rom_array[25296] = 32'hFFFFFFF1;
    // rom_array[25297] = 32'hFFFFFFF1;
    // rom_array[25298] = 32'hFFFFFFF1;
    // rom_array[25299] = 32'hFFFFFFF1;
    // rom_array[25300] = 32'hFFFFFFF1;
    // rom_array[25301] = 32'hFFFFFFF1;
    // rom_array[25302] = 32'hFFFFFFF1;
    // rom_array[25303] = 32'hFFFFFFF1;
    // rom_array[25304] = 32'hFFFFFFF1;
    // rom_array[25305] = 32'hFFFFFFF1;
    // rom_array[25306] = 32'hFFFFFFF1;
    // rom_array[25307] = 32'hFFFFFFF1;
    // rom_array[25308] = 32'hFFFFFFF1;
    // rom_array[25309] = 32'hFFFFFFF1;
    // rom_array[25310] = 32'hFFFFFFF1;
    // rom_array[25311] = 32'hFFFFFFF1;
    // rom_array[25312] = 32'hFFFFFFF1;
    // rom_array[25313] = 32'hFFFFFFF1;
    // rom_array[25314] = 32'hFFFFFFF1;
    // rom_array[25315] = 32'hFFFFFFF1;
    // rom_array[25316] = 32'hFFFFFFF1;
    // rom_array[25317] = 32'hFFFFFFF1;
    // rom_array[25318] = 32'hFFFFFFF1;
    // rom_array[25319] = 32'hFFFFFFF1;
    // rom_array[25320] = 32'hFFFFFFF1;
    // rom_array[25321] = 32'hFFFFFFF1;
    // rom_array[25322] = 32'hFFFFFFF1;
    // rom_array[25323] = 32'hFFFFFFF1;
    // rom_array[25324] = 32'hFFFFFFF1;
    // rom_array[25325] = 32'hFFFFFFF1;
    // rom_array[25326] = 32'hFFFFFFF1;
    // rom_array[25327] = 32'hFFFFFFF1;
    // rom_array[25328] = 32'hFFFFFFF1;
    // rom_array[25329] = 32'hFFFFFFF1;
    // rom_array[25330] = 32'hFFFFFFF1;
    // rom_array[25331] = 32'hFFFFFFF1;
    // rom_array[25332] = 32'hFFFFFFF1;
    // rom_array[25333] = 32'hFFFFFFF1;
    // rom_array[25334] = 32'hFFFFFFF1;
    // rom_array[25335] = 32'hFFFFFFF1;
    // rom_array[25336] = 32'hFFFFFFF1;
    // rom_array[25337] = 32'hFFFFFFF1;
    // rom_array[25338] = 32'hFFFFFFF1;
    // rom_array[25339] = 32'hFFFFFFF1;
    // rom_array[25340] = 32'hFFFFFFF1;
    // rom_array[25341] = 32'hFFFFFFF1;
    // rom_array[25342] = 32'hFFFFFFF1;
    // rom_array[25343] = 32'hFFFFFFF1;
    // rom_array[25344] = 32'hFFFFFFF1;
    // rom_array[25345] = 32'hFFFFFFF1;
    // rom_array[25346] = 32'hFFFFFFF1;
    // rom_array[25347] = 32'hFFFFFFF1;
    // rom_array[25348] = 32'hFFFFFFF1;
    // rom_array[25349] = 32'hFFFFFFF1;
    // rom_array[25350] = 32'hFFFFFFF1;
    // rom_array[25351] = 32'hFFFFFFF1;
    // rom_array[25352] = 32'hFFFFFFF1;
    // rom_array[25353] = 32'hFFFFFFF0;
    // rom_array[25354] = 32'hFFFFFFF0;
    // rom_array[25355] = 32'hFFFFFFF0;
    // rom_array[25356] = 32'hFFFFFFF0;
    // rom_array[25357] = 32'hFFFFFFF0;
    // rom_array[25358] = 32'hFFFFFFF0;
    // rom_array[25359] = 32'hFFFFFFF1;
    // rom_array[25360] = 32'hFFFFFFF1;
    // rom_array[25361] = 32'hFFFFFFF0;
    // rom_array[25362] = 32'hFFFFFFF0;
    // rom_array[25363] = 32'hFFFFFFF0;
    // rom_array[25364] = 32'hFFFFFFF0;
    // rom_array[25365] = 32'hFFFFFFF0;
    // rom_array[25366] = 32'hFFFFFFF0;
    // rom_array[25367] = 32'hFFFFFFF1;
    // rom_array[25368] = 32'hFFFFFFF1;
    // rom_array[25369] = 32'hFFFFFFF0;
    // rom_array[25370] = 32'hFFFFFFF0;
    // rom_array[25371] = 32'hFFFFFFF0;
    // rom_array[25372] = 32'hFFFFFFF0;
    // rom_array[25373] = 32'hFFFFFFF1;
    // rom_array[25374] = 32'hFFFFFFF1;
    // rom_array[25375] = 32'hFFFFFFF1;
    // rom_array[25376] = 32'hFFFFFFF1;
    // rom_array[25377] = 32'hFFFFFFF0;
    // rom_array[25378] = 32'hFFFFFFF0;
    // rom_array[25379] = 32'hFFFFFFF0;
    // rom_array[25380] = 32'hFFFFFFF0;
    // rom_array[25381] = 32'hFFFFFFF1;
    // rom_array[25382] = 32'hFFFFFFF1;
    // rom_array[25383] = 32'hFFFFFFF1;
    // rom_array[25384] = 32'hFFFFFFF1;
    // rom_array[25385] = 32'hFFFFFFF0;
    // rom_array[25386] = 32'hFFFFFFF0;
    // rom_array[25387] = 32'hFFFFFFF1;
    // rom_array[25388] = 32'hFFFFFFF1;
    // rom_array[25389] = 32'hFFFFFFF0;
    // rom_array[25390] = 32'hFFFFFFF0;
    // rom_array[25391] = 32'hFFFFFFF1;
    // rom_array[25392] = 32'hFFFFFFF1;
    // rom_array[25393] = 32'hFFFFFFF0;
    // rom_array[25394] = 32'hFFFFFFF0;
    // rom_array[25395] = 32'hFFFFFFF1;
    // rom_array[25396] = 32'hFFFFFFF1;
    // rom_array[25397] = 32'hFFFFFFF0;
    // rom_array[25398] = 32'hFFFFFFF0;
    // rom_array[25399] = 32'hFFFFFFF1;
    // rom_array[25400] = 32'hFFFFFFF1;
    // rom_array[25401] = 32'hFFFFFFF0;
    // rom_array[25402] = 32'hFFFFFFF0;
    // rom_array[25403] = 32'hFFFFFFF1;
    // rom_array[25404] = 32'hFFFFFFF1;
    // rom_array[25405] = 32'hFFFFFFF0;
    // rom_array[25406] = 32'hFFFFFFF0;
    // rom_array[25407] = 32'hFFFFFFF1;
    // rom_array[25408] = 32'hFFFFFFF1;
    // rom_array[25409] = 32'hFFFFFFF0;
    // rom_array[25410] = 32'hFFFFFFF0;
    // rom_array[25411] = 32'hFFFFFFF1;
    // rom_array[25412] = 32'hFFFFFFF1;
    // rom_array[25413] = 32'hFFFFFFF0;
    // rom_array[25414] = 32'hFFFFFFF0;
    // rom_array[25415] = 32'hFFFFFFF1;
    // rom_array[25416] = 32'hFFFFFFF1;
    // rom_array[25417] = 32'hFFFFFFF0;
    // rom_array[25418] = 32'hFFFFFFF0;
    // rom_array[25419] = 32'hFFFFFFF0;
    // rom_array[25420] = 32'hFFFFFFF0;
    // rom_array[25421] = 32'hFFFFFFF1;
    // rom_array[25422] = 32'hFFFFFFF1;
    // rom_array[25423] = 32'hFFFFFFF1;
    // rom_array[25424] = 32'hFFFFFFF1;
    // rom_array[25425] = 32'hFFFFFFF0;
    // rom_array[25426] = 32'hFFFFFFF0;
    // rom_array[25427] = 32'hFFFFFFF0;
    // rom_array[25428] = 32'hFFFFFFF0;
    // rom_array[25429] = 32'hFFFFFFF1;
    // rom_array[25430] = 32'hFFFFFFF1;
    // rom_array[25431] = 32'hFFFFFFF1;
    // rom_array[25432] = 32'hFFFFFFF1;
    // rom_array[25433] = 32'hFFFFFFF0;
    // rom_array[25434] = 32'hFFFFFFF0;
    // rom_array[25435] = 32'hFFFFFFF0;
    // rom_array[25436] = 32'hFFFFFFF0;
    // rom_array[25437] = 32'hFFFFFFF1;
    // rom_array[25438] = 32'hFFFFFFF1;
    // rom_array[25439] = 32'hFFFFFFF1;
    // rom_array[25440] = 32'hFFFFFFF1;
    // rom_array[25441] = 32'hFFFFFFF0;
    // rom_array[25442] = 32'hFFFFFFF0;
    // rom_array[25443] = 32'hFFFFFFF0;
    // rom_array[25444] = 32'hFFFFFFF0;
    // rom_array[25445] = 32'hFFFFFFF1;
    // rom_array[25446] = 32'hFFFFFFF1;
    // rom_array[25447] = 32'hFFFFFFF1;
    // rom_array[25448] = 32'hFFFFFFF1;
    // rom_array[25449] = 32'hFFFFFFF0;
    // rom_array[25450] = 32'hFFFFFFF0;
    // rom_array[25451] = 32'hFFFFFFF0;
    // rom_array[25452] = 32'hFFFFFFF0;
    // rom_array[25453] = 32'hFFFFFFF1;
    // rom_array[25454] = 32'hFFFFFFF1;
    // rom_array[25455] = 32'hFFFFFFF1;
    // rom_array[25456] = 32'hFFFFFFF1;
    // rom_array[25457] = 32'hFFFFFFF0;
    // rom_array[25458] = 32'hFFFFFFF0;
    // rom_array[25459] = 32'hFFFFFFF0;
    // rom_array[25460] = 32'hFFFFFFF0;
    // rom_array[25461] = 32'hFFFFFFF1;
    // rom_array[25462] = 32'hFFFFFFF1;
    // rom_array[25463] = 32'hFFFFFFF1;
    // rom_array[25464] = 32'hFFFFFFF1;
    // rom_array[25465] = 32'hFFFFFFF1;
    // rom_array[25466] = 32'hFFFFFFF1;
    // rom_array[25467] = 32'hFFFFFFF1;
    // rom_array[25468] = 32'hFFFFFFF1;
    // rom_array[25469] = 32'hFFFFFFF1;
    // rom_array[25470] = 32'hFFFFFFF1;
    // rom_array[25471] = 32'hFFFFFFF1;
    // rom_array[25472] = 32'hFFFFFFF1;
    // rom_array[25473] = 32'hFFFFFFF1;
    // rom_array[25474] = 32'hFFFFFFF1;
    // rom_array[25475] = 32'hFFFFFFF1;
    // rom_array[25476] = 32'hFFFFFFF1;
    // rom_array[25477] = 32'hFFFFFFF1;
    // rom_array[25478] = 32'hFFFFFFF1;
    // rom_array[25479] = 32'hFFFFFFF1;
    // rom_array[25480] = 32'hFFFFFFF1;
    // rom_array[25481] = 32'hFFFFFFF1;
    // rom_array[25482] = 32'hFFFFFFF1;
    // rom_array[25483] = 32'hFFFFFFF1;
    // rom_array[25484] = 32'hFFFFFFF1;
    // rom_array[25485] = 32'hFFFFFFF1;
    // rom_array[25486] = 32'hFFFFFFF1;
    // rom_array[25487] = 32'hFFFFFFF1;
    // rom_array[25488] = 32'hFFFFFFF1;
    // rom_array[25489] = 32'hFFFFFFF1;
    // rom_array[25490] = 32'hFFFFFFF1;
    // rom_array[25491] = 32'hFFFFFFF1;
    // rom_array[25492] = 32'hFFFFFFF1;
    // rom_array[25493] = 32'hFFFFFFF1;
    // rom_array[25494] = 32'hFFFFFFF1;
    // rom_array[25495] = 32'hFFFFFFF1;
    // rom_array[25496] = 32'hFFFFFFF1;
    // rom_array[25497] = 32'hFFFFFFF0;
    // rom_array[25498] = 32'hFFFFFFF0;
    // rom_array[25499] = 32'hFFFFFFF0;
    // rom_array[25500] = 32'hFFFFFFF0;
    // rom_array[25501] = 32'hFFFFFFF1;
    // rom_array[25502] = 32'hFFFFFFF1;
    // rom_array[25503] = 32'hFFFFFFF1;
    // rom_array[25504] = 32'hFFFFFFF1;
    // rom_array[25505] = 32'hFFFFFFF0;
    // rom_array[25506] = 32'hFFFFFFF0;
    // rom_array[25507] = 32'hFFFFFFF0;
    // rom_array[25508] = 32'hFFFFFFF0;
    // rom_array[25509] = 32'hFFFFFFF1;
    // rom_array[25510] = 32'hFFFFFFF1;
    // rom_array[25511] = 32'hFFFFFFF1;
    // rom_array[25512] = 32'hFFFFFFF1;
    // rom_array[25513] = 32'hFFFFFFF0;
    // rom_array[25514] = 32'hFFFFFFF0;
    // rom_array[25515] = 32'hFFFFFFF0;
    // rom_array[25516] = 32'hFFFFFFF0;
    // rom_array[25517] = 32'hFFFFFFF1;
    // rom_array[25518] = 32'hFFFFFFF1;
    // rom_array[25519] = 32'hFFFFFFF1;
    // rom_array[25520] = 32'hFFFFFFF1;
    // rom_array[25521] = 32'hFFFFFFF0;
    // rom_array[25522] = 32'hFFFFFFF0;
    // rom_array[25523] = 32'hFFFFFFF0;
    // rom_array[25524] = 32'hFFFFFFF0;
    // rom_array[25525] = 32'hFFFFFFF1;
    // rom_array[25526] = 32'hFFFFFFF1;
    // rom_array[25527] = 32'hFFFFFFF1;
    // rom_array[25528] = 32'hFFFFFFF1;
    // rom_array[25529] = 32'hFFFFFFF0;
    // rom_array[25530] = 32'hFFFFFFF0;
    // rom_array[25531] = 32'hFFFFFFF0;
    // rom_array[25532] = 32'hFFFFFFF0;
    // rom_array[25533] = 32'hFFFFFFF1;
    // rom_array[25534] = 32'hFFFFFFF1;
    // rom_array[25535] = 32'hFFFFFFF1;
    // rom_array[25536] = 32'hFFFFFFF1;
    // rom_array[25537] = 32'hFFFFFFF0;
    // rom_array[25538] = 32'hFFFFFFF0;
    // rom_array[25539] = 32'hFFFFFFF0;
    // rom_array[25540] = 32'hFFFFFFF0;
    // rom_array[25541] = 32'hFFFFFFF1;
    // rom_array[25542] = 32'hFFFFFFF1;
    // rom_array[25543] = 32'hFFFFFFF1;
    // rom_array[25544] = 32'hFFFFFFF1;
    // rom_array[25545] = 32'hFFFFFFF0;
    // rom_array[25546] = 32'hFFFFFFF0;
    // rom_array[25547] = 32'hFFFFFFF0;
    // rom_array[25548] = 32'hFFFFFFF0;
    // rom_array[25549] = 32'hFFFFFFF1;
    // rom_array[25550] = 32'hFFFFFFF1;
    // rom_array[25551] = 32'hFFFFFFF1;
    // rom_array[25552] = 32'hFFFFFFF1;
    // rom_array[25553] = 32'hFFFFFFF0;
    // rom_array[25554] = 32'hFFFFFFF0;
    // rom_array[25555] = 32'hFFFFFFF0;
    // rom_array[25556] = 32'hFFFFFFF0;
    // rom_array[25557] = 32'hFFFFFFF1;
    // rom_array[25558] = 32'hFFFFFFF1;
    // rom_array[25559] = 32'hFFFFFFF1;
    // rom_array[25560] = 32'hFFFFFFF1;
    // rom_array[25561] = 32'hFFFFFFF0;
    // rom_array[25562] = 32'hFFFFFFF0;
    // rom_array[25563] = 32'hFFFFFFF1;
    // rom_array[25564] = 32'hFFFFFFF1;
    // rom_array[25565] = 32'hFFFFFFF0;
    // rom_array[25566] = 32'hFFFFFFF0;
    // rom_array[25567] = 32'hFFFFFFF1;
    // rom_array[25568] = 32'hFFFFFFF1;
    // rom_array[25569] = 32'hFFFFFFF0;
    // rom_array[25570] = 32'hFFFFFFF0;
    // rom_array[25571] = 32'hFFFFFFF1;
    // rom_array[25572] = 32'hFFFFFFF1;
    // rom_array[25573] = 32'hFFFFFFF0;
    // rom_array[25574] = 32'hFFFFFFF0;
    // rom_array[25575] = 32'hFFFFFFF1;
    // rom_array[25576] = 32'hFFFFFFF1;
    // rom_array[25577] = 32'hFFFFFFF0;
    // rom_array[25578] = 32'hFFFFFFF0;
    // rom_array[25579] = 32'hFFFFFFF1;
    // rom_array[25580] = 32'hFFFFFFF1;
    // rom_array[25581] = 32'hFFFFFFF0;
    // rom_array[25582] = 32'hFFFFFFF0;
    // rom_array[25583] = 32'hFFFFFFF1;
    // rom_array[25584] = 32'hFFFFFFF1;
    // rom_array[25585] = 32'hFFFFFFF0;
    // rom_array[25586] = 32'hFFFFFFF0;
    // rom_array[25587] = 32'hFFFFFFF1;
    // rom_array[25588] = 32'hFFFFFFF1;
    // rom_array[25589] = 32'hFFFFFFF0;
    // rom_array[25590] = 32'hFFFFFFF0;
    // rom_array[25591] = 32'hFFFFFFF1;
    // rom_array[25592] = 32'hFFFFFFF1;
    // rom_array[25593] = 32'hFFFFFFF0;
    // rom_array[25594] = 32'hFFFFFFF0;
    // rom_array[25595] = 32'hFFFFFFF0;
    // rom_array[25596] = 32'hFFFFFFF0;
    // rom_array[25597] = 32'hFFFFFFF1;
    // rom_array[25598] = 32'hFFFFFFF1;
    // rom_array[25599] = 32'hFFFFFFF1;
    // rom_array[25600] = 32'hFFFFFFF1;
    // rom_array[25601] = 32'hFFFFFFF0;
    // rom_array[25602] = 32'hFFFFFFF0;
    // rom_array[25603] = 32'hFFFFFFF0;
    // rom_array[25604] = 32'hFFFFFFF0;
    // rom_array[25605] = 32'hFFFFFFF1;
    // rom_array[25606] = 32'hFFFFFFF1;
    // rom_array[25607] = 32'hFFFFFFF1;
    // rom_array[25608] = 32'hFFFFFFF1;
    // rom_array[25609] = 32'hFFFFFFF0;
    // rom_array[25610] = 32'hFFFFFFF0;
    // rom_array[25611] = 32'hFFFFFFF0;
    // rom_array[25612] = 32'hFFFFFFF0;
    // rom_array[25613] = 32'hFFFFFFF1;
    // rom_array[25614] = 32'hFFFFFFF1;
    // rom_array[25615] = 32'hFFFFFFF1;
    // rom_array[25616] = 32'hFFFFFFF1;
    // rom_array[25617] = 32'hFFFFFFF0;
    // rom_array[25618] = 32'hFFFFFFF0;
    // rom_array[25619] = 32'hFFFFFFF0;
    // rom_array[25620] = 32'hFFFFFFF0;
    // rom_array[25621] = 32'hFFFFFFF1;
    // rom_array[25622] = 32'hFFFFFFF1;
    // rom_array[25623] = 32'hFFFFFFF1;
    // rom_array[25624] = 32'hFFFFFFF1;
    // rom_array[25625] = 32'hFFFFFFF0;
    // rom_array[25626] = 32'hFFFFFFF0;
    // rom_array[25627] = 32'hFFFFFFF1;
    // rom_array[25628] = 32'hFFFFFFF1;
    // rom_array[25629] = 32'hFFFFFFF1;
    // rom_array[25630] = 32'hFFFFFFF1;
    // rom_array[25631] = 32'hFFFFFFF1;
    // rom_array[25632] = 32'hFFFFFFF1;
    // rom_array[25633] = 32'hFFFFFFF0;
    // rom_array[25634] = 32'hFFFFFFF0;
    // rom_array[25635] = 32'hFFFFFFF1;
    // rom_array[25636] = 32'hFFFFFFF1;
    // rom_array[25637] = 32'hFFFFFFF1;
    // rom_array[25638] = 32'hFFFFFFF1;
    // rom_array[25639] = 32'hFFFFFFF1;
    // rom_array[25640] = 32'hFFFFFFF1;
    // rom_array[25641] = 32'hFFFFFFF1;
    // rom_array[25642] = 32'hFFFFFFF1;
    // rom_array[25643] = 32'hFFFFFFF1;
    // rom_array[25644] = 32'hFFFFFFF1;
    // rom_array[25645] = 32'hFFFFFFF1;
    // rom_array[25646] = 32'hFFFFFFF1;
    // rom_array[25647] = 32'hFFFFFFF1;
    // rom_array[25648] = 32'hFFFFFFF1;
    // rom_array[25649] = 32'hFFFFFFF1;
    // rom_array[25650] = 32'hFFFFFFF1;
    // rom_array[25651] = 32'hFFFFFFF1;
    // rom_array[25652] = 32'hFFFFFFF1;
    // rom_array[25653] = 32'hFFFFFFF1;
    // rom_array[25654] = 32'hFFFFFFF1;
    // rom_array[25655] = 32'hFFFFFFF1;
    // rom_array[25656] = 32'hFFFFFFF1;
    // rom_array[25657] = 32'hFFFFFFF1;
    // rom_array[25658] = 32'hFFFFFFF1;
    // rom_array[25659] = 32'hFFFFFFF1;
    // rom_array[25660] = 32'hFFFFFFF1;
    // rom_array[25661] = 32'hFFFFFFF0;
    // rom_array[25662] = 32'hFFFFFFF0;
    // rom_array[25663] = 32'hFFFFFFF0;
    // rom_array[25664] = 32'hFFFFFFF0;
    // rom_array[25665] = 32'hFFFFFFF1;
    // rom_array[25666] = 32'hFFFFFFF1;
    // rom_array[25667] = 32'hFFFFFFF1;
    // rom_array[25668] = 32'hFFFFFFF1;
    // rom_array[25669] = 32'hFFFFFFF0;
    // rom_array[25670] = 32'hFFFFFFF0;
    // rom_array[25671] = 32'hFFFFFFF0;
    // rom_array[25672] = 32'hFFFFFFF0;
    // rom_array[25673] = 32'hFFFFFFF1;
    // rom_array[25674] = 32'hFFFFFFF1;
    // rom_array[25675] = 32'hFFFFFFF1;
    // rom_array[25676] = 32'hFFFFFFF1;
    // rom_array[25677] = 32'hFFFFFFF0;
    // rom_array[25678] = 32'hFFFFFFF0;
    // rom_array[25679] = 32'hFFFFFFF0;
    // rom_array[25680] = 32'hFFFFFFF0;
    // rom_array[25681] = 32'hFFFFFFF1;
    // rom_array[25682] = 32'hFFFFFFF1;
    // rom_array[25683] = 32'hFFFFFFF1;
    // rom_array[25684] = 32'hFFFFFFF1;
    // rom_array[25685] = 32'hFFFFFFF0;
    // rom_array[25686] = 32'hFFFFFFF0;
    // rom_array[25687] = 32'hFFFFFFF0;
    // rom_array[25688] = 32'hFFFFFFF0;
    // rom_array[25689] = 32'hFFFFFFF1;
    // rom_array[25690] = 32'hFFFFFFF1;
    // rom_array[25691] = 32'hFFFFFFF1;
    // rom_array[25692] = 32'hFFFFFFF1;
    // rom_array[25693] = 32'hFFFFFFF0;
    // rom_array[25694] = 32'hFFFFFFF0;
    // rom_array[25695] = 32'hFFFFFFF0;
    // rom_array[25696] = 32'hFFFFFFF0;
    // rom_array[25697] = 32'hFFFFFFF1;
    // rom_array[25698] = 32'hFFFFFFF1;
    // rom_array[25699] = 32'hFFFFFFF1;
    // rom_array[25700] = 32'hFFFFFFF1;
    // rom_array[25701] = 32'hFFFFFFF0;
    // rom_array[25702] = 32'hFFFFFFF0;
    // rom_array[25703] = 32'hFFFFFFF0;
    // rom_array[25704] = 32'hFFFFFFF0;
    // rom_array[25705] = 32'hFFFFFFF1;
    // rom_array[25706] = 32'hFFFFFFF1;
    // rom_array[25707] = 32'hFFFFFFF1;
    // rom_array[25708] = 32'hFFFFFFF1;
    // rom_array[25709] = 32'hFFFFFFF0;
    // rom_array[25710] = 32'hFFFFFFF0;
    // rom_array[25711] = 32'hFFFFFFF0;
    // rom_array[25712] = 32'hFFFFFFF0;
    // rom_array[25713] = 32'hFFFFFFF1;
    // rom_array[25714] = 32'hFFFFFFF1;
    // rom_array[25715] = 32'hFFFFFFF1;
    // rom_array[25716] = 32'hFFFFFFF1;
    // rom_array[25717] = 32'hFFFFFFF0;
    // rom_array[25718] = 32'hFFFFFFF0;
    // rom_array[25719] = 32'hFFFFFFF0;
    // rom_array[25720] = 32'hFFFFFFF0;
    // rom_array[25721] = 32'hFFFFFFF1;
    // rom_array[25722] = 32'hFFFFFFF1;
    // rom_array[25723] = 32'hFFFFFFF1;
    // rom_array[25724] = 32'hFFFFFFF1;
    // rom_array[25725] = 32'hFFFFFFF1;
    // rom_array[25726] = 32'hFFFFFFF1;
    // rom_array[25727] = 32'hFFFFFFF1;
    // rom_array[25728] = 32'hFFFFFFF1;
    // rom_array[25729] = 32'hFFFFFFF1;
    // rom_array[25730] = 32'hFFFFFFF1;
    // rom_array[25731] = 32'hFFFFFFF1;
    // rom_array[25732] = 32'hFFFFFFF1;
    // rom_array[25733] = 32'hFFFFFFF1;
    // rom_array[25734] = 32'hFFFFFFF1;
    // rom_array[25735] = 32'hFFFFFFF1;
    // rom_array[25736] = 32'hFFFFFFF1;
    // rom_array[25737] = 32'hFFFFFFF1;
    // rom_array[25738] = 32'hFFFFFFF1;
    // rom_array[25739] = 32'hFFFFFFF1;
    // rom_array[25740] = 32'hFFFFFFF1;
    // rom_array[25741] = 32'hFFFFFFF1;
    // rom_array[25742] = 32'hFFFFFFF1;
    // rom_array[25743] = 32'hFFFFFFF1;
    // rom_array[25744] = 32'hFFFFFFF1;
    // rom_array[25745] = 32'hFFFFFFF1;
    // rom_array[25746] = 32'hFFFFFFF1;
    // rom_array[25747] = 32'hFFFFFFF1;
    // rom_array[25748] = 32'hFFFFFFF1;
    // rom_array[25749] = 32'hFFFFFFF1;
    // rom_array[25750] = 32'hFFFFFFF1;
    // rom_array[25751] = 32'hFFFFFFF1;
    // rom_array[25752] = 32'hFFFFFFF1;
    // rom_array[25753] = 32'hFFFFFFF1;
    // rom_array[25754] = 32'hFFFFFFF1;
    // rom_array[25755] = 32'hFFFFFFF1;
    // rom_array[25756] = 32'hFFFFFFF1;
    // rom_array[25757] = 32'hFFFFFFF0;
    // rom_array[25758] = 32'hFFFFFFF0;
    // rom_array[25759] = 32'hFFFFFFF0;
    // rom_array[25760] = 32'hFFFFFFF0;
    // rom_array[25761] = 32'hFFFFFFF1;
    // rom_array[25762] = 32'hFFFFFFF1;
    // rom_array[25763] = 32'hFFFFFFF1;
    // rom_array[25764] = 32'hFFFFFFF1;
    // rom_array[25765] = 32'hFFFFFFF0;
    // rom_array[25766] = 32'hFFFFFFF0;
    // rom_array[25767] = 32'hFFFFFFF0;
    // rom_array[25768] = 32'hFFFFFFF0;
    // rom_array[25769] = 32'hFFFFFFF1;
    // rom_array[25770] = 32'hFFFFFFF1;
    // rom_array[25771] = 32'hFFFFFFF1;
    // rom_array[25772] = 32'hFFFFFFF1;
    // rom_array[25773] = 32'hFFFFFFF0;
    // rom_array[25774] = 32'hFFFFFFF0;
    // rom_array[25775] = 32'hFFFFFFF0;
    // rom_array[25776] = 32'hFFFFFFF0;
    // rom_array[25777] = 32'hFFFFFFF1;
    // rom_array[25778] = 32'hFFFFFFF1;
    // rom_array[25779] = 32'hFFFFFFF1;
    // rom_array[25780] = 32'hFFFFFFF1;
    // rom_array[25781] = 32'hFFFFFFF0;
    // rom_array[25782] = 32'hFFFFFFF0;
    // rom_array[25783] = 32'hFFFFFFF0;
    // rom_array[25784] = 32'hFFFFFFF0;
    // rom_array[25785] = 32'hFFFFFFF1;
    // rom_array[25786] = 32'hFFFFFFF1;
    // rom_array[25787] = 32'hFFFFFFF1;
    // rom_array[25788] = 32'hFFFFFFF1;
    // rom_array[25789] = 32'hFFFFFFF0;
    // rom_array[25790] = 32'hFFFFFFF0;
    // rom_array[25791] = 32'hFFFFFFF1;
    // rom_array[25792] = 32'hFFFFFFF1;
    // rom_array[25793] = 32'hFFFFFFF1;
    // rom_array[25794] = 32'hFFFFFFF1;
    // rom_array[25795] = 32'hFFFFFFF1;
    // rom_array[25796] = 32'hFFFFFFF1;
    // rom_array[25797] = 32'hFFFFFFF0;
    // rom_array[25798] = 32'hFFFFFFF0;
    // rom_array[25799] = 32'hFFFFFFF1;
    // rom_array[25800] = 32'hFFFFFFF1;
    // rom_array[25801] = 32'hFFFFFFF0;
    // rom_array[25802] = 32'hFFFFFFF0;
    // rom_array[25803] = 32'hFFFFFFF1;
    // rom_array[25804] = 32'hFFFFFFF1;
    // rom_array[25805] = 32'hFFFFFFF0;
    // rom_array[25806] = 32'hFFFFFFF0;
    // rom_array[25807] = 32'hFFFFFFF1;
    // rom_array[25808] = 32'hFFFFFFF1;
    // rom_array[25809] = 32'hFFFFFFF0;
    // rom_array[25810] = 32'hFFFFFFF0;
    // rom_array[25811] = 32'hFFFFFFF1;
    // rom_array[25812] = 32'hFFFFFFF1;
    // rom_array[25813] = 32'hFFFFFFF0;
    // rom_array[25814] = 32'hFFFFFFF0;
    // rom_array[25815] = 32'hFFFFFFF1;
    // rom_array[25816] = 32'hFFFFFFF1;
    // rom_array[25817] = 32'hFFFFFFF1;
    // rom_array[25818] = 32'hFFFFFFF1;
    // rom_array[25819] = 32'hFFFFFFF1;
    // rom_array[25820] = 32'hFFFFFFF1;
    // rom_array[25821] = 32'hFFFFFFF1;
    // rom_array[25822] = 32'hFFFFFFF1;
    // rom_array[25823] = 32'hFFFFFFF1;
    // rom_array[25824] = 32'hFFFFFFF1;
    // rom_array[25825] = 32'hFFFFFFF1;
    // rom_array[25826] = 32'hFFFFFFF1;
    // rom_array[25827] = 32'hFFFFFFF1;
    // rom_array[25828] = 32'hFFFFFFF1;
    // rom_array[25829] = 32'hFFFFFFF1;
    // rom_array[25830] = 32'hFFFFFFF1;
    // rom_array[25831] = 32'hFFFFFFF1;
    // rom_array[25832] = 32'hFFFFFFF1;
    // rom_array[25833] = 32'hFFFFFFF1;
    // rom_array[25834] = 32'hFFFFFFF1;
    // rom_array[25835] = 32'hFFFFFFF1;
    // rom_array[25836] = 32'hFFFFFFF1;
    // rom_array[25837] = 32'hFFFFFFF1;
    // rom_array[25838] = 32'hFFFFFFF1;
    // rom_array[25839] = 32'hFFFFFFF1;
    // rom_array[25840] = 32'hFFFFFFF1;
    // rom_array[25841] = 32'hFFFFFFF1;
    // rom_array[25842] = 32'hFFFFFFF1;
    // rom_array[25843] = 32'hFFFFFFF1;
    // rom_array[25844] = 32'hFFFFFFF1;
    // rom_array[25845] = 32'hFFFFFFF1;
    // rom_array[25846] = 32'hFFFFFFF1;
    // rom_array[25847] = 32'hFFFFFFF1;
    // rom_array[25848] = 32'hFFFFFFF1;
    // rom_array[25849] = 32'hFFFFFFF1;
    // rom_array[25850] = 32'hFFFFFFF1;
    // rom_array[25851] = 32'hFFFFFFF1;
    // rom_array[25852] = 32'hFFFFFFF1;
    // rom_array[25853] = 32'hFFFFFFF1;
    // rom_array[25854] = 32'hFFFFFFF1;
    // rom_array[25855] = 32'hFFFFFFF1;
    // rom_array[25856] = 32'hFFFFFFF1;
    // rom_array[25857] = 32'hFFFFFFF1;
    // rom_array[25858] = 32'hFFFFFFF1;
    // rom_array[25859] = 32'hFFFFFFF1;
    // rom_array[25860] = 32'hFFFFFFF1;
    // rom_array[25861] = 32'hFFFFFFF1;
    // rom_array[25862] = 32'hFFFFFFF1;
    // rom_array[25863] = 32'hFFFFFFF1;
    // rom_array[25864] = 32'hFFFFFFF1;
    // rom_array[25865] = 32'hFFFFFFF1;
    // rom_array[25866] = 32'hFFFFFFF1;
    // rom_array[25867] = 32'hFFFFFFF1;
    // rom_array[25868] = 32'hFFFFFFF1;
    // rom_array[25869] = 32'hFFFFFFF1;
    // rom_array[25870] = 32'hFFFFFFF1;
    // rom_array[25871] = 32'hFFFFFFF1;
    // rom_array[25872] = 32'hFFFFFFF1;
    // rom_array[25873] = 32'hFFFFFFF1;
    // rom_array[25874] = 32'hFFFFFFF1;
    // rom_array[25875] = 32'hFFFFFFF1;
    // rom_array[25876] = 32'hFFFFFFF1;
    // rom_array[25877] = 32'hFFFFFFF1;
    // rom_array[25878] = 32'hFFFFFFF1;
    // rom_array[25879] = 32'hFFFFFFF1;
    // rom_array[25880] = 32'hFFFFFFF1;
    // rom_array[25881] = 32'hFFFFFFF1;
    // rom_array[25882] = 32'hFFFFFFF1;
    // rom_array[25883] = 32'hFFFFFFF1;
    // rom_array[25884] = 32'hFFFFFFF1;
    // rom_array[25885] = 32'hFFFFFFF1;
    // rom_array[25886] = 32'hFFFFFFF1;
    // rom_array[25887] = 32'hFFFFFFF1;
    // rom_array[25888] = 32'hFFFFFFF1;
    // rom_array[25889] = 32'hFFFFFFF1;
    // rom_array[25890] = 32'hFFFFFFF1;
    // rom_array[25891] = 32'hFFFFFFF1;
    // rom_array[25892] = 32'hFFFFFFF1;
    // rom_array[25893] = 32'hFFFFFFF1;
    // rom_array[25894] = 32'hFFFFFFF1;
    // rom_array[25895] = 32'hFFFFFFF1;
    // rom_array[25896] = 32'hFFFFFFF1;
    // rom_array[25897] = 32'hFFFFFFF1;
    // rom_array[25898] = 32'hFFFFFFF1;
    // rom_array[25899] = 32'hFFFFFFF1;
    // rom_array[25900] = 32'hFFFFFFF1;
    // rom_array[25901] = 32'hFFFFFFF1;
    // rom_array[25902] = 32'hFFFFFFF1;
    // rom_array[25903] = 32'hFFFFFFF1;
    // rom_array[25904] = 32'hFFFFFFF1;
    // rom_array[25905] = 32'hFFFFFFF1;
    // rom_array[25906] = 32'hFFFFFFF1;
    // rom_array[25907] = 32'hFFFFFFF1;
    // rom_array[25908] = 32'hFFFFFFF1;
    // rom_array[25909] = 32'hFFFFFFF1;
    // rom_array[25910] = 32'hFFFFFFF1;
    // rom_array[25911] = 32'hFFFFFFF1;
    // rom_array[25912] = 32'hFFFFFFF1;
    // rom_array[25913] = 32'hFFFFFFF1;
    // rom_array[25914] = 32'hFFFFFFF1;
    // rom_array[25915] = 32'hFFFFFFF1;
    // rom_array[25916] = 32'hFFFFFFF1;
    // rom_array[25917] = 32'hFFFFFFF1;
    // rom_array[25918] = 32'hFFFFFFF1;
    // rom_array[25919] = 32'hFFFFFFF1;
    // rom_array[25920] = 32'hFFFFFFF1;
    // rom_array[25921] = 32'hFFFFFFF1;
    // rom_array[25922] = 32'hFFFFFFF1;
    // rom_array[25923] = 32'hFFFFFFF1;
    // rom_array[25924] = 32'hFFFFFFF1;
    // rom_array[25925] = 32'hFFFFFFF1;
    // rom_array[25926] = 32'hFFFFFFF1;
    // rom_array[25927] = 32'hFFFFFFF1;
    // rom_array[25928] = 32'hFFFFFFF1;
    // rom_array[25929] = 32'hFFFFFFF1;
    // rom_array[25930] = 32'hFFFFFFF1;
    // rom_array[25931] = 32'hFFFFFFF1;
    // rom_array[25932] = 32'hFFFFFFF1;
    // rom_array[25933] = 32'hFFFFFFF1;
    // rom_array[25934] = 32'hFFFFFFF1;
    // rom_array[25935] = 32'hFFFFFFF1;
    // rom_array[25936] = 32'hFFFFFFF1;
    // rom_array[25937] = 32'hFFFFFFF1;
    // rom_array[25938] = 32'hFFFFFFF1;
    // rom_array[25939] = 32'hFFFFFFF1;
    // rom_array[25940] = 32'hFFFFFFF1;
    // rom_array[25941] = 32'hFFFFFFF1;
    // rom_array[25942] = 32'hFFFFFFF1;
    // rom_array[25943] = 32'hFFFFFFF1;
    // rom_array[25944] = 32'hFFFFFFF1;
    // rom_array[25945] = 32'hFFFFFFF0;
    // rom_array[25946] = 32'hFFFFFFF0;
    // rom_array[25947] = 32'hFFFFFFF1;
    // rom_array[25948] = 32'hFFFFFFF1;
    // rom_array[25949] = 32'hFFFFFFF0;
    // rom_array[25950] = 32'hFFFFFFF0;
    // rom_array[25951] = 32'hFFFFFFF1;
    // rom_array[25952] = 32'hFFFFFFF1;
    // rom_array[25953] = 32'hFFFFFFF0;
    // rom_array[25954] = 32'hFFFFFFF0;
    // rom_array[25955] = 32'hFFFFFFF1;
    // rom_array[25956] = 32'hFFFFFFF1;
    // rom_array[25957] = 32'hFFFFFFF0;
    // rom_array[25958] = 32'hFFFFFFF0;
    // rom_array[25959] = 32'hFFFFFFF1;
    // rom_array[25960] = 32'hFFFFFFF1;
    // rom_array[25961] = 32'hFFFFFFF0;
    // rom_array[25962] = 32'hFFFFFFF0;
    // rom_array[25963] = 32'hFFFFFFF1;
    // rom_array[25964] = 32'hFFFFFFF1;
    // rom_array[25965] = 32'hFFFFFFF0;
    // rom_array[25966] = 32'hFFFFFFF0;
    // rom_array[25967] = 32'hFFFFFFF1;
    // rom_array[25968] = 32'hFFFFFFF1;
    // rom_array[25969] = 32'hFFFFFFF0;
    // rom_array[25970] = 32'hFFFFFFF0;
    // rom_array[25971] = 32'hFFFFFFF1;
    // rom_array[25972] = 32'hFFFFFFF1;
    // rom_array[25973] = 32'hFFFFFFF0;
    // rom_array[25974] = 32'hFFFFFFF0;
    // rom_array[25975] = 32'hFFFFFFF1;
    // rom_array[25976] = 32'hFFFFFFF1;
    // rom_array[25977] = 32'hFFFFFFF0;
    // rom_array[25978] = 32'hFFFFFFF0;
    // rom_array[25979] = 32'hFFFFFFF1;
    // rom_array[25980] = 32'hFFFFFFF1;
    // rom_array[25981] = 32'hFFFFFFF0;
    // rom_array[25982] = 32'hFFFFFFF0;
    // rom_array[25983] = 32'hFFFFFFF1;
    // rom_array[25984] = 32'hFFFFFFF1;
    // rom_array[25985] = 32'hFFFFFFF0;
    // rom_array[25986] = 32'hFFFFFFF0;
    // rom_array[25987] = 32'hFFFFFFF1;
    // rom_array[25988] = 32'hFFFFFFF1;
    // rom_array[25989] = 32'hFFFFFFF0;
    // rom_array[25990] = 32'hFFFFFFF0;
    // rom_array[25991] = 32'hFFFFFFF1;
    // rom_array[25992] = 32'hFFFFFFF1;
    // rom_array[25993] = 32'hFFFFFFF0;
    // rom_array[25994] = 32'hFFFFFFF0;
    // rom_array[25995] = 32'hFFFFFFF1;
    // rom_array[25996] = 32'hFFFFFFF1;
    // rom_array[25997] = 32'hFFFFFFF0;
    // rom_array[25998] = 32'hFFFFFFF0;
    // rom_array[25999] = 32'hFFFFFFF0;
    // rom_array[26000] = 32'hFFFFFFF0;
    // rom_array[26001] = 32'hFFFFFFF0;
    // rom_array[26002] = 32'hFFFFFFF0;
    // rom_array[26003] = 32'hFFFFFFF1;
    // rom_array[26004] = 32'hFFFFFFF1;
    // rom_array[26005] = 32'hFFFFFFF0;
    // rom_array[26006] = 32'hFFFFFFF0;
    // rom_array[26007] = 32'hFFFFFFF0;
    // rom_array[26008] = 32'hFFFFFFF0;
    // rom_array[26009] = 32'hFFFFFFF1;
    // rom_array[26010] = 32'hFFFFFFF1;
    // rom_array[26011] = 32'hFFFFFFF1;
    // rom_array[26012] = 32'hFFFFFFF1;
    // rom_array[26013] = 32'hFFFFFFF0;
    // rom_array[26014] = 32'hFFFFFFF0;
    // rom_array[26015] = 32'hFFFFFFF0;
    // rom_array[26016] = 32'hFFFFFFF0;
    // rom_array[26017] = 32'hFFFFFFF1;
    // rom_array[26018] = 32'hFFFFFFF1;
    // rom_array[26019] = 32'hFFFFFFF1;
    // rom_array[26020] = 32'hFFFFFFF1;
    // rom_array[26021] = 32'hFFFFFFF0;
    // rom_array[26022] = 32'hFFFFFFF0;
    // rom_array[26023] = 32'hFFFFFFF0;
    // rom_array[26024] = 32'hFFFFFFF0;
    // rom_array[26025] = 32'hFFFFFFF1;
    // rom_array[26026] = 32'hFFFFFFF1;
    // rom_array[26027] = 32'hFFFFFFF1;
    // rom_array[26028] = 32'hFFFFFFF1;
    // rom_array[26029] = 32'hFFFFFFF1;
    // rom_array[26030] = 32'hFFFFFFF1;
    // rom_array[26031] = 32'hFFFFFFF1;
    // rom_array[26032] = 32'hFFFFFFF1;
    // rom_array[26033] = 32'hFFFFFFF1;
    // rom_array[26034] = 32'hFFFFFFF1;
    // rom_array[26035] = 32'hFFFFFFF1;
    // rom_array[26036] = 32'hFFFFFFF1;
    // rom_array[26037] = 32'hFFFFFFF1;
    // rom_array[26038] = 32'hFFFFFFF1;
    // rom_array[26039] = 32'hFFFFFFF1;
    // rom_array[26040] = 32'hFFFFFFF1;
    // rom_array[26041] = 32'hFFFFFFF1;
    // rom_array[26042] = 32'hFFFFFFF1;
    // rom_array[26043] = 32'hFFFFFFF1;
    // rom_array[26044] = 32'hFFFFFFF1;
    // rom_array[26045] = 32'hFFFFFFF1;
    // rom_array[26046] = 32'hFFFFFFF1;
    // rom_array[26047] = 32'hFFFFFFF1;
    // rom_array[26048] = 32'hFFFFFFF1;
    // rom_array[26049] = 32'hFFFFFFF1;
    // rom_array[26050] = 32'hFFFFFFF1;
    // rom_array[26051] = 32'hFFFFFFF1;
    // rom_array[26052] = 32'hFFFFFFF1;
    // rom_array[26053] = 32'hFFFFFFF1;
    // rom_array[26054] = 32'hFFFFFFF1;
    // rom_array[26055] = 32'hFFFFFFF1;
    // rom_array[26056] = 32'hFFFFFFF1;
    // rom_array[26057] = 32'hFFFFFFF1;
    // rom_array[26058] = 32'hFFFFFFF1;
    // rom_array[26059] = 32'hFFFFFFF1;
    // rom_array[26060] = 32'hFFFFFFF1;
    // rom_array[26061] = 32'hFFFFFFF0;
    // rom_array[26062] = 32'hFFFFFFF0;
    // rom_array[26063] = 32'hFFFFFFF0;
    // rom_array[26064] = 32'hFFFFFFF0;
    // rom_array[26065] = 32'hFFFFFFF1;
    // rom_array[26066] = 32'hFFFFFFF1;
    // rom_array[26067] = 32'hFFFFFFF1;
    // rom_array[26068] = 32'hFFFFFFF1;
    // rom_array[26069] = 32'hFFFFFFF0;
    // rom_array[26070] = 32'hFFFFFFF0;
    // rom_array[26071] = 32'hFFFFFFF0;
    // rom_array[26072] = 32'hFFFFFFF0;
    // rom_array[26073] = 32'hFFFFFFF1;
    // rom_array[26074] = 32'hFFFFFFF1;
    // rom_array[26075] = 32'hFFFFFFF1;
    // rom_array[26076] = 32'hFFFFFFF1;
    // rom_array[26077] = 32'hFFFFFFF0;
    // rom_array[26078] = 32'hFFFFFFF0;
    // rom_array[26079] = 32'hFFFFFFF0;
    // rom_array[26080] = 32'hFFFFFFF0;
    // rom_array[26081] = 32'hFFFFFFF1;
    // rom_array[26082] = 32'hFFFFFFF1;
    // rom_array[26083] = 32'hFFFFFFF1;
    // rom_array[26084] = 32'hFFFFFFF1;
    // rom_array[26085] = 32'hFFFFFFF0;
    // rom_array[26086] = 32'hFFFFFFF0;
    // rom_array[26087] = 32'hFFFFFFF0;
    // rom_array[26088] = 32'hFFFFFFF0;
    // rom_array[26089] = 32'hFFFFFFF1;
    // rom_array[26090] = 32'hFFFFFFF1;
    // rom_array[26091] = 32'hFFFFFFF1;
    // rom_array[26092] = 32'hFFFFFFF1;
    // rom_array[26093] = 32'hFFFFFFF1;
    // rom_array[26094] = 32'hFFFFFFF1;
    // rom_array[26095] = 32'hFFFFFFF1;
    // rom_array[26096] = 32'hFFFFFFF1;
    // rom_array[26097] = 32'hFFFFFFF1;
    // rom_array[26098] = 32'hFFFFFFF1;
    // rom_array[26099] = 32'hFFFFFFF1;
    // rom_array[26100] = 32'hFFFFFFF1;
    // rom_array[26101] = 32'hFFFFFFF1;
    // rom_array[26102] = 32'hFFFFFFF1;
    // rom_array[26103] = 32'hFFFFFFF1;
    // rom_array[26104] = 32'hFFFFFFF1;
    // rom_array[26105] = 32'hFFFFFFF1;
    // rom_array[26106] = 32'hFFFFFFF1;
    // rom_array[26107] = 32'hFFFFFFF1;
    // rom_array[26108] = 32'hFFFFFFF1;
    // rom_array[26109] = 32'hFFFFFFF0;
    // rom_array[26110] = 32'hFFFFFFF0;
    // rom_array[26111] = 32'hFFFFFFF0;
    // rom_array[26112] = 32'hFFFFFFF0;
    // rom_array[26113] = 32'hFFFFFFF1;
    // rom_array[26114] = 32'hFFFFFFF1;
    // rom_array[26115] = 32'hFFFFFFF1;
    // rom_array[26116] = 32'hFFFFFFF1;
    // rom_array[26117] = 32'hFFFFFFF0;
    // rom_array[26118] = 32'hFFFFFFF0;
    // rom_array[26119] = 32'hFFFFFFF0;
    // rom_array[26120] = 32'hFFFFFFF0;
    // rom_array[26121] = 32'hFFFFFFF0;
    // rom_array[26122] = 32'hFFFFFFF0;
    // rom_array[26123] = 32'hFFFFFFF0;
    // rom_array[26124] = 32'hFFFFFFF0;
    // rom_array[26125] = 32'hFFFFFFF1;
    // rom_array[26126] = 32'hFFFFFFF1;
    // rom_array[26127] = 32'hFFFFFFF1;
    // rom_array[26128] = 32'hFFFFFFF1;
    // rom_array[26129] = 32'hFFFFFFF0;
    // rom_array[26130] = 32'hFFFFFFF0;
    // rom_array[26131] = 32'hFFFFFFF0;
    // rom_array[26132] = 32'hFFFFFFF0;
    // rom_array[26133] = 32'hFFFFFFF1;
    // rom_array[26134] = 32'hFFFFFFF1;
    // rom_array[26135] = 32'hFFFFFFF1;
    // rom_array[26136] = 32'hFFFFFFF1;
    // rom_array[26137] = 32'hFFFFFFF0;
    // rom_array[26138] = 32'hFFFFFFF0;
    // rom_array[26139] = 32'hFFFFFFF0;
    // rom_array[26140] = 32'hFFFFFFF0;
    // rom_array[26141] = 32'hFFFFFFF1;
    // rom_array[26142] = 32'hFFFFFFF1;
    // rom_array[26143] = 32'hFFFFFFF1;
    // rom_array[26144] = 32'hFFFFFFF1;
    // rom_array[26145] = 32'hFFFFFFF0;
    // rom_array[26146] = 32'hFFFFFFF0;
    // rom_array[26147] = 32'hFFFFFFF0;
    // rom_array[26148] = 32'hFFFFFFF0;
    // rom_array[26149] = 32'hFFFFFFF1;
    // rom_array[26150] = 32'hFFFFFFF1;
    // rom_array[26151] = 32'hFFFFFFF1;
    // rom_array[26152] = 32'hFFFFFFF1;
    // rom_array[26153] = 32'hFFFFFFF1;
    // rom_array[26154] = 32'hFFFFFFF1;
    // rom_array[26155] = 32'hFFFFFFF1;
    // rom_array[26156] = 32'hFFFFFFF1;
    // rom_array[26157] = 32'hFFFFFFF1;
    // rom_array[26158] = 32'hFFFFFFF1;
    // rom_array[26159] = 32'hFFFFFFF1;
    // rom_array[26160] = 32'hFFFFFFF1;
    // rom_array[26161] = 32'hFFFFFFF1;
    // rom_array[26162] = 32'hFFFFFFF1;
    // rom_array[26163] = 32'hFFFFFFF1;
    // rom_array[26164] = 32'hFFFFFFF1;
    // rom_array[26165] = 32'hFFFFFFF1;
    // rom_array[26166] = 32'hFFFFFFF1;
    // rom_array[26167] = 32'hFFFFFFF1;
    // rom_array[26168] = 32'hFFFFFFF1;
    // rom_array[26169] = 32'hFFFFFFF1;
    // rom_array[26170] = 32'hFFFFFFF1;
    // rom_array[26171] = 32'hFFFFFFF1;
    // rom_array[26172] = 32'hFFFFFFF1;
    // rom_array[26173] = 32'hFFFFFFF1;
    // rom_array[26174] = 32'hFFFFFFF1;
    // rom_array[26175] = 32'hFFFFFFF1;
    // rom_array[26176] = 32'hFFFFFFF1;
    // rom_array[26177] = 32'hFFFFFFF1;
    // rom_array[26178] = 32'hFFFFFFF1;
    // rom_array[26179] = 32'hFFFFFFF1;
    // rom_array[26180] = 32'hFFFFFFF1;
    // rom_array[26181] = 32'hFFFFFFF1;
    // rom_array[26182] = 32'hFFFFFFF1;
    // rom_array[26183] = 32'hFFFFFFF1;
    // rom_array[26184] = 32'hFFFFFFF1;
    // rom_array[26185] = 32'hFFFFFFF0;
    // rom_array[26186] = 32'hFFFFFFF0;
    // rom_array[26187] = 32'hFFFFFFF0;
    // rom_array[26188] = 32'hFFFFFFF0;
    // rom_array[26189] = 32'hFFFFFFF1;
    // rom_array[26190] = 32'hFFFFFFF1;
    // rom_array[26191] = 32'hFFFFFFF1;
    // rom_array[26192] = 32'hFFFFFFF1;
    // rom_array[26193] = 32'hFFFFFFF0;
    // rom_array[26194] = 32'hFFFFFFF0;
    // rom_array[26195] = 32'hFFFFFFF0;
    // rom_array[26196] = 32'hFFFFFFF0;
    // rom_array[26197] = 32'hFFFFFFF1;
    // rom_array[26198] = 32'hFFFFFFF1;
    // rom_array[26199] = 32'hFFFFFFF1;
    // rom_array[26200] = 32'hFFFFFFF1;
    // rom_array[26201] = 32'hFFFFFFF0;
    // rom_array[26202] = 32'hFFFFFFF0;
    // rom_array[26203] = 32'hFFFFFFF0;
    // rom_array[26204] = 32'hFFFFFFF0;
    // rom_array[26205] = 32'hFFFFFFF1;
    // rom_array[26206] = 32'hFFFFFFF1;
    // rom_array[26207] = 32'hFFFFFFF1;
    // rom_array[26208] = 32'hFFFFFFF1;
    // rom_array[26209] = 32'hFFFFFFF0;
    // rom_array[26210] = 32'hFFFFFFF0;
    // rom_array[26211] = 32'hFFFFFFF0;
    // rom_array[26212] = 32'hFFFFFFF0;
    // rom_array[26213] = 32'hFFFFFFF1;
    // rom_array[26214] = 32'hFFFFFFF1;
    // rom_array[26215] = 32'hFFFFFFF1;
    // rom_array[26216] = 32'hFFFFFFF1;
    // rom_array[26217] = 32'hFFFFFFF1;
    // rom_array[26218] = 32'hFFFFFFF1;
    // rom_array[26219] = 32'hFFFFFFF1;
    // rom_array[26220] = 32'hFFFFFFF1;
    // rom_array[26221] = 32'hFFFFFFF1;
    // rom_array[26222] = 32'hFFFFFFF1;
    // rom_array[26223] = 32'hFFFFFFF1;
    // rom_array[26224] = 32'hFFFFFFF1;
    // rom_array[26225] = 32'hFFFFFFF1;
    // rom_array[26226] = 32'hFFFFFFF1;
    // rom_array[26227] = 32'hFFFFFFF1;
    // rom_array[26228] = 32'hFFFFFFF1;
    // rom_array[26229] = 32'hFFFFFFF1;
    // rom_array[26230] = 32'hFFFFFFF1;
    // rom_array[26231] = 32'hFFFFFFF1;
    // rom_array[26232] = 32'hFFFFFFF1;
    // rom_array[26233] = 32'hFFFFFFF1;
    // rom_array[26234] = 32'hFFFFFFF1;
    // rom_array[26235] = 32'hFFFFFFF1;
    // rom_array[26236] = 32'hFFFFFFF1;
    // rom_array[26237] = 32'hFFFFFFF1;
    // rom_array[26238] = 32'hFFFFFFF1;
    // rom_array[26239] = 32'hFFFFFFF1;
    // rom_array[26240] = 32'hFFFFFFF1;
    // rom_array[26241] = 32'hFFFFFFF1;
    // rom_array[26242] = 32'hFFFFFFF1;
    // rom_array[26243] = 32'hFFFFFFF1;
    // rom_array[26244] = 32'hFFFFFFF1;
    // rom_array[26245] = 32'hFFFFFFF1;
    // rom_array[26246] = 32'hFFFFFFF1;
    // rom_array[26247] = 32'hFFFFFFF1;
    // rom_array[26248] = 32'hFFFFFFF1;
    // rom_array[26249] = 32'hFFFFFFF0;
    // rom_array[26250] = 32'hFFFFFFF0;
    // rom_array[26251] = 32'hFFFFFFF0;
    // rom_array[26252] = 32'hFFFFFFF0;
    // rom_array[26253] = 32'hFFFFFFF1;
    // rom_array[26254] = 32'hFFFFFFF1;
    // rom_array[26255] = 32'hFFFFFFF1;
    // rom_array[26256] = 32'hFFFFFFF1;
    // rom_array[26257] = 32'hFFFFFFF0;
    // rom_array[26258] = 32'hFFFFFFF0;
    // rom_array[26259] = 32'hFFFFFFF0;
    // rom_array[26260] = 32'hFFFFFFF0;
    // rom_array[26261] = 32'hFFFFFFF1;
    // rom_array[26262] = 32'hFFFFFFF1;
    // rom_array[26263] = 32'hFFFFFFF1;
    // rom_array[26264] = 32'hFFFFFFF1;
    // rom_array[26265] = 32'hFFFFFFF0;
    // rom_array[26266] = 32'hFFFFFFF0;
    // rom_array[26267] = 32'hFFFFFFF0;
    // rom_array[26268] = 32'hFFFFFFF0;
    // rom_array[26269] = 32'hFFFFFFF1;
    // rom_array[26270] = 32'hFFFFFFF1;
    // rom_array[26271] = 32'hFFFFFFF1;
    // rom_array[26272] = 32'hFFFFFFF1;
    // rom_array[26273] = 32'hFFFFFFF0;
    // rom_array[26274] = 32'hFFFFFFF0;
    // rom_array[26275] = 32'hFFFFFFF0;
    // rom_array[26276] = 32'hFFFFFFF0;
    // rom_array[26277] = 32'hFFFFFFF1;
    // rom_array[26278] = 32'hFFFFFFF1;
    // rom_array[26279] = 32'hFFFFFFF1;
    // rom_array[26280] = 32'hFFFFFFF1;
    // rom_array[26281] = 32'hFFFFFFF1;
    // rom_array[26282] = 32'hFFFFFFF1;
    // rom_array[26283] = 32'hFFFFFFF1;
    // rom_array[26284] = 32'hFFFFFFF1;
    // rom_array[26285] = 32'hFFFFFFF1;
    // rom_array[26286] = 32'hFFFFFFF1;
    // rom_array[26287] = 32'hFFFFFFF1;
    // rom_array[26288] = 32'hFFFFFFF1;
    // rom_array[26289] = 32'hFFFFFFF1;
    // rom_array[26290] = 32'hFFFFFFF1;
    // rom_array[26291] = 32'hFFFFFFF1;
    // rom_array[26292] = 32'hFFFFFFF1;
    // rom_array[26293] = 32'hFFFFFFF1;
    // rom_array[26294] = 32'hFFFFFFF1;
    // rom_array[26295] = 32'hFFFFFFF1;
    // rom_array[26296] = 32'hFFFFFFF1;
    // rom_array[26297] = 32'hFFFFFFF1;
    // rom_array[26298] = 32'hFFFFFFF1;
    // rom_array[26299] = 32'hFFFFFFF1;
    // rom_array[26300] = 32'hFFFFFFF1;
    // rom_array[26301] = 32'hFFFFFFF1;
    // rom_array[26302] = 32'hFFFFFFF1;
    // rom_array[26303] = 32'hFFFFFFF1;
    // rom_array[26304] = 32'hFFFFFFF1;
    // rom_array[26305] = 32'hFFFFFFF1;
    // rom_array[26306] = 32'hFFFFFFF1;
    // rom_array[26307] = 32'hFFFFFFF1;
    // rom_array[26308] = 32'hFFFFFFF1;
    // rom_array[26309] = 32'hFFFFFFF1;
    // rom_array[26310] = 32'hFFFFFFF1;
    // rom_array[26311] = 32'hFFFFFFF1;
    // rom_array[26312] = 32'hFFFFFFF1;
    // rom_array[26313] = 32'hFFFFFFF0;
    // rom_array[26314] = 32'hFFFFFFF0;
    // rom_array[26315] = 32'hFFFFFFF0;
    // rom_array[26316] = 32'hFFFFFFF0;
    // rom_array[26317] = 32'hFFFFFFF1;
    // rom_array[26318] = 32'hFFFFFFF1;
    // rom_array[26319] = 32'hFFFFFFF1;
    // rom_array[26320] = 32'hFFFFFFF1;
    // rom_array[26321] = 32'hFFFFFFF0;
    // rom_array[26322] = 32'hFFFFFFF0;
    // rom_array[26323] = 32'hFFFFFFF0;
    // rom_array[26324] = 32'hFFFFFFF0;
    // rom_array[26325] = 32'hFFFFFFF1;
    // rom_array[26326] = 32'hFFFFFFF1;
    // rom_array[26327] = 32'hFFFFFFF1;
    // rom_array[26328] = 32'hFFFFFFF1;
    // rom_array[26329] = 32'hFFFFFFF0;
    // rom_array[26330] = 32'hFFFFFFF0;
    // rom_array[26331] = 32'hFFFFFFF0;
    // rom_array[26332] = 32'hFFFFFFF0;
    // rom_array[26333] = 32'hFFFFFFF1;
    // rom_array[26334] = 32'hFFFFFFF1;
    // rom_array[26335] = 32'hFFFFFFF1;
    // rom_array[26336] = 32'hFFFFFFF1;
    // rom_array[26337] = 32'hFFFFFFF0;
    // rom_array[26338] = 32'hFFFFFFF0;
    // rom_array[26339] = 32'hFFFFFFF0;
    // rom_array[26340] = 32'hFFFFFFF0;
    // rom_array[26341] = 32'hFFFFFFF1;
    // rom_array[26342] = 32'hFFFFFFF1;
    // rom_array[26343] = 32'hFFFFFFF1;
    // rom_array[26344] = 32'hFFFFFFF1;
    // rom_array[26345] = 32'hFFFFFFF1;
    // rom_array[26346] = 32'hFFFFFFF1;
    // rom_array[26347] = 32'hFFFFFFF1;
    // rom_array[26348] = 32'hFFFFFFF1;
    // rom_array[26349] = 32'hFFFFFFF1;
    // rom_array[26350] = 32'hFFFFFFF1;
    // rom_array[26351] = 32'hFFFFFFF1;
    // rom_array[26352] = 32'hFFFFFFF1;
    // rom_array[26353] = 32'hFFFFFFF1;
    // rom_array[26354] = 32'hFFFFFFF1;
    // rom_array[26355] = 32'hFFFFFFF1;
    // rom_array[26356] = 32'hFFFFFFF1;
    // rom_array[26357] = 32'hFFFFFFF1;
    // rom_array[26358] = 32'hFFFFFFF1;
    // rom_array[26359] = 32'hFFFFFFF1;
    // rom_array[26360] = 32'hFFFFFFF1;
    // rom_array[26361] = 32'hFFFFFFF1;
    // rom_array[26362] = 32'hFFFFFFF1;
    // rom_array[26363] = 32'hFFFFFFF1;
    // rom_array[26364] = 32'hFFFFFFF1;
    // rom_array[26365] = 32'hFFFFFFF1;
    // rom_array[26366] = 32'hFFFFFFF1;
    // rom_array[26367] = 32'hFFFFFFF1;
    // rom_array[26368] = 32'hFFFFFFF1;
    // rom_array[26369] = 32'hFFFFFFF1;
    // rom_array[26370] = 32'hFFFFFFF1;
    // rom_array[26371] = 32'hFFFFFFF1;
    // rom_array[26372] = 32'hFFFFFFF1;
    // rom_array[26373] = 32'hFFFFFFF1;
    // rom_array[26374] = 32'hFFFFFFF1;
    // rom_array[26375] = 32'hFFFFFFF1;
    // rom_array[26376] = 32'hFFFFFFF1;
    // rom_array[26377] = 32'hFFFFFFF0;
    // rom_array[26378] = 32'hFFFFFFF0;
    // rom_array[26379] = 32'hFFFFFFF0;
    // rom_array[26380] = 32'hFFFFFFF0;
    // rom_array[26381] = 32'hFFFFFFF1;
    // rom_array[26382] = 32'hFFFFFFF1;
    // rom_array[26383] = 32'hFFFFFFF1;
    // rom_array[26384] = 32'hFFFFFFF1;
    // rom_array[26385] = 32'hFFFFFFF0;
    // rom_array[26386] = 32'hFFFFFFF0;
    // rom_array[26387] = 32'hFFFFFFF0;
    // rom_array[26388] = 32'hFFFFFFF0;
    // rom_array[26389] = 32'hFFFFFFF1;
    // rom_array[26390] = 32'hFFFFFFF1;
    // rom_array[26391] = 32'hFFFFFFF1;
    // rom_array[26392] = 32'hFFFFFFF1;
    // rom_array[26393] = 32'hFFFFFFF0;
    // rom_array[26394] = 32'hFFFFFFF0;
    // rom_array[26395] = 32'hFFFFFFF0;
    // rom_array[26396] = 32'hFFFFFFF0;
    // rom_array[26397] = 32'hFFFFFFF1;
    // rom_array[26398] = 32'hFFFFFFF1;
    // rom_array[26399] = 32'hFFFFFFF1;
    // rom_array[26400] = 32'hFFFFFFF1;
    // rom_array[26401] = 32'hFFFFFFF0;
    // rom_array[26402] = 32'hFFFFFFF0;
    // rom_array[26403] = 32'hFFFFFFF0;
    // rom_array[26404] = 32'hFFFFFFF0;
    // rom_array[26405] = 32'hFFFFFFF1;
    // rom_array[26406] = 32'hFFFFFFF1;
    // rom_array[26407] = 32'hFFFFFFF1;
    // rom_array[26408] = 32'hFFFFFFF1;
    // rom_array[26409] = 32'hFFFFFFF1;
    // rom_array[26410] = 32'hFFFFFFF1;
    // rom_array[26411] = 32'hFFFFFFF1;
    // rom_array[26412] = 32'hFFFFFFF1;
    // rom_array[26413] = 32'hFFFFFFF1;
    // rom_array[26414] = 32'hFFFFFFF1;
    // rom_array[26415] = 32'hFFFFFFF1;
    // rom_array[26416] = 32'hFFFFFFF1;
    // rom_array[26417] = 32'hFFFFFFF1;
    // rom_array[26418] = 32'hFFFFFFF1;
    // rom_array[26419] = 32'hFFFFFFF1;
    // rom_array[26420] = 32'hFFFFFFF1;
    // rom_array[26421] = 32'hFFFFFFF1;
    // rom_array[26422] = 32'hFFFFFFF1;
    // rom_array[26423] = 32'hFFFFFFF1;
    // rom_array[26424] = 32'hFFFFFFF1;
    // rom_array[26425] = 32'hFFFFFFF1;
    // rom_array[26426] = 32'hFFFFFFF1;
    // rom_array[26427] = 32'hFFFFFFF1;
    // rom_array[26428] = 32'hFFFFFFF1;
    // rom_array[26429] = 32'hFFFFFFF1;
    // rom_array[26430] = 32'hFFFFFFF1;
    // rom_array[26431] = 32'hFFFFFFF1;
    // rom_array[26432] = 32'hFFFFFFF1;
    // rom_array[26433] = 32'hFFFFFFF1;
    // rom_array[26434] = 32'hFFFFFFF1;
    // rom_array[26435] = 32'hFFFFFFF1;
    // rom_array[26436] = 32'hFFFFFFF1;
    // rom_array[26437] = 32'hFFFFFFF1;
    // rom_array[26438] = 32'hFFFFFFF1;
    // rom_array[26439] = 32'hFFFFFFF1;
    // rom_array[26440] = 32'hFFFFFFF1;
    // rom_array[26441] = 32'hFFFFFFF0;
    // rom_array[26442] = 32'hFFFFFFF0;
    // rom_array[26443] = 32'hFFFFFFF0;
    // rom_array[26444] = 32'hFFFFFFF0;
    // rom_array[26445] = 32'hFFFFFFF1;
    // rom_array[26446] = 32'hFFFFFFF1;
    // rom_array[26447] = 32'hFFFFFFF1;
    // rom_array[26448] = 32'hFFFFFFF1;
    // rom_array[26449] = 32'hFFFFFFF0;
    // rom_array[26450] = 32'hFFFFFFF0;
    // rom_array[26451] = 32'hFFFFFFF0;
    // rom_array[26452] = 32'hFFFFFFF0;
    // rom_array[26453] = 32'hFFFFFFF1;
    // rom_array[26454] = 32'hFFFFFFF1;
    // rom_array[26455] = 32'hFFFFFFF1;
    // rom_array[26456] = 32'hFFFFFFF1;
    // rom_array[26457] = 32'hFFFFFFF1;
    // rom_array[26458] = 32'hFFFFFFF1;
    // rom_array[26459] = 32'hFFFFFFF1;
    // rom_array[26460] = 32'hFFFFFFF1;
    // rom_array[26461] = 32'hFFFFFFF1;
    // rom_array[26462] = 32'hFFFFFFF1;
    // rom_array[26463] = 32'hFFFFFFF1;
    // rom_array[26464] = 32'hFFFFFFF1;
    // rom_array[26465] = 32'hFFFFFFF1;
    // rom_array[26466] = 32'hFFFFFFF1;
    // rom_array[26467] = 32'hFFFFFFF1;
    // rom_array[26468] = 32'hFFFFFFF1;
    // rom_array[26469] = 32'hFFFFFFF1;
    // rom_array[26470] = 32'hFFFFFFF1;
    // rom_array[26471] = 32'hFFFFFFF1;
    // rom_array[26472] = 32'hFFFFFFF1;
    // rom_array[26473] = 32'hFFFFFFF1;
    // rom_array[26474] = 32'hFFFFFFF1;
    // rom_array[26475] = 32'hFFFFFFF0;
    // rom_array[26476] = 32'hFFFFFFF0;
    // rom_array[26477] = 32'hFFFFFFF1;
    // rom_array[26478] = 32'hFFFFFFF1;
    // rom_array[26479] = 32'hFFFFFFF0;
    // rom_array[26480] = 32'hFFFFFFF0;
    // rom_array[26481] = 32'hFFFFFFF1;
    // rom_array[26482] = 32'hFFFFFFF1;
    // rom_array[26483] = 32'hFFFFFFF0;
    // rom_array[26484] = 32'hFFFFFFF0;
    // rom_array[26485] = 32'hFFFFFFF1;
    // rom_array[26486] = 32'hFFFFFFF1;
    // rom_array[26487] = 32'hFFFFFFF0;
    // rom_array[26488] = 32'hFFFFFFF0;
    // rom_array[26489] = 32'hFFFFFFF1;
    // rom_array[26490] = 32'hFFFFFFF1;
    // rom_array[26491] = 32'hFFFFFFF1;
    // rom_array[26492] = 32'hFFFFFFF1;
    // rom_array[26493] = 32'hFFFFFFF0;
    // rom_array[26494] = 32'hFFFFFFF0;
    // rom_array[26495] = 32'hFFFFFFF0;
    // rom_array[26496] = 32'hFFFFFFF0;
    // rom_array[26497] = 32'hFFFFFFF1;
    // rom_array[26498] = 32'hFFFFFFF1;
    // rom_array[26499] = 32'hFFFFFFF1;
    // rom_array[26500] = 32'hFFFFFFF1;
    // rom_array[26501] = 32'hFFFFFFF0;
    // rom_array[26502] = 32'hFFFFFFF0;
    // rom_array[26503] = 32'hFFFFFFF0;
    // rom_array[26504] = 32'hFFFFFFF0;
    // rom_array[26505] = 32'hFFFFFFF1;
    // rom_array[26506] = 32'hFFFFFFF1;
    // rom_array[26507] = 32'hFFFFFFF1;
    // rom_array[26508] = 32'hFFFFFFF1;
    // rom_array[26509] = 32'hFFFFFFF0;
    // rom_array[26510] = 32'hFFFFFFF0;
    // rom_array[26511] = 32'hFFFFFFF0;
    // rom_array[26512] = 32'hFFFFFFF0;
    // rom_array[26513] = 32'hFFFFFFF1;
    // rom_array[26514] = 32'hFFFFFFF1;
    // rom_array[26515] = 32'hFFFFFFF1;
    // rom_array[26516] = 32'hFFFFFFF1;
    // rom_array[26517] = 32'hFFFFFFF0;
    // rom_array[26518] = 32'hFFFFFFF0;
    // rom_array[26519] = 32'hFFFFFFF0;
    // rom_array[26520] = 32'hFFFFFFF0;
    // rom_array[26521] = 32'hFFFFFFF1;
    // rom_array[26522] = 32'hFFFFFFF1;
    // rom_array[26523] = 32'hFFFFFFF1;
    // rom_array[26524] = 32'hFFFFFFF1;
    // rom_array[26525] = 32'hFFFFFFF0;
    // rom_array[26526] = 32'hFFFFFFF0;
    // rom_array[26527] = 32'hFFFFFFF0;
    // rom_array[26528] = 32'hFFFFFFF0;
    // rom_array[26529] = 32'hFFFFFFF1;
    // rom_array[26530] = 32'hFFFFFFF1;
    // rom_array[26531] = 32'hFFFFFFF1;
    // rom_array[26532] = 32'hFFFFFFF1;
    // rom_array[26533] = 32'hFFFFFFF0;
    // rom_array[26534] = 32'hFFFFFFF0;
    // rom_array[26535] = 32'hFFFFFFF0;
    // rom_array[26536] = 32'hFFFFFFF0;
    // rom_array[26537] = 32'hFFFFFFF1;
    // rom_array[26538] = 32'hFFFFFFF1;
    // rom_array[26539] = 32'hFFFFFFF1;
    // rom_array[26540] = 32'hFFFFFFF1;
    // rom_array[26541] = 32'hFFFFFFF0;
    // rom_array[26542] = 32'hFFFFFFF0;
    // rom_array[26543] = 32'hFFFFFFF0;
    // rom_array[26544] = 32'hFFFFFFF0;
    // rom_array[26545] = 32'hFFFFFFF1;
    // rom_array[26546] = 32'hFFFFFFF1;
    // rom_array[26547] = 32'hFFFFFFF1;
    // rom_array[26548] = 32'hFFFFFFF1;
    // rom_array[26549] = 32'hFFFFFFF0;
    // rom_array[26550] = 32'hFFFFFFF0;
    // rom_array[26551] = 32'hFFFFFFF0;
    // rom_array[26552] = 32'hFFFFFFF0;
    // rom_array[26553] = 32'hFFFFFFF1;
    // rom_array[26554] = 32'hFFFFFFF1;
    // rom_array[26555] = 32'hFFFFFFF1;
    // rom_array[26556] = 32'hFFFFFFF1;
    // rom_array[26557] = 32'hFFFFFFF0;
    // rom_array[26558] = 32'hFFFFFFF0;
    // rom_array[26559] = 32'hFFFFFFF0;
    // rom_array[26560] = 32'hFFFFFFF0;
    // rom_array[26561] = 32'hFFFFFFF1;
    // rom_array[26562] = 32'hFFFFFFF1;
    // rom_array[26563] = 32'hFFFFFFF1;
    // rom_array[26564] = 32'hFFFFFFF1;
    // rom_array[26565] = 32'hFFFFFFF0;
    // rom_array[26566] = 32'hFFFFFFF0;
    // rom_array[26567] = 32'hFFFFFFF0;
    // rom_array[26568] = 32'hFFFFFFF0;
    // rom_array[26569] = 32'hFFFFFFF1;
    // rom_array[26570] = 32'hFFFFFFF1;
    // rom_array[26571] = 32'hFFFFFFF1;
    // rom_array[26572] = 32'hFFFFFFF1;
    // rom_array[26573] = 32'hFFFFFFF0;
    // rom_array[26574] = 32'hFFFFFFF0;
    // rom_array[26575] = 32'hFFFFFFF0;
    // rom_array[26576] = 32'hFFFFFFF0;
    // rom_array[26577] = 32'hFFFFFFF1;
    // rom_array[26578] = 32'hFFFFFFF1;
    // rom_array[26579] = 32'hFFFFFFF1;
    // rom_array[26580] = 32'hFFFFFFF1;
    // rom_array[26581] = 32'hFFFFFFF0;
    // rom_array[26582] = 32'hFFFFFFF0;
    // rom_array[26583] = 32'hFFFFFFF0;
    // rom_array[26584] = 32'hFFFFFFF0;
    // rom_array[26585] = 32'hFFFFFFF1;
    // rom_array[26586] = 32'hFFFFFFF1;
    // rom_array[26587] = 32'hFFFFFFF1;
    // rom_array[26588] = 32'hFFFFFFF1;
    // rom_array[26589] = 32'hFFFFFFF0;
    // rom_array[26590] = 32'hFFFFFFF0;
    // rom_array[26591] = 32'hFFFFFFF0;
    // rom_array[26592] = 32'hFFFFFFF0;
    // rom_array[26593] = 32'hFFFFFFF1;
    // rom_array[26594] = 32'hFFFFFFF1;
    // rom_array[26595] = 32'hFFFFFFF1;
    // rom_array[26596] = 32'hFFFFFFF1;
    // rom_array[26597] = 32'hFFFFFFF0;
    // rom_array[26598] = 32'hFFFFFFF0;
    // rom_array[26599] = 32'hFFFFFFF0;
    // rom_array[26600] = 32'hFFFFFFF0;
    // rom_array[26601] = 32'hFFFFFFF1;
    // rom_array[26602] = 32'hFFFFFFF1;
    // rom_array[26603] = 32'hFFFFFFF1;
    // rom_array[26604] = 32'hFFFFFFF1;
    // rom_array[26605] = 32'hFFFFFFF0;
    // rom_array[26606] = 32'hFFFFFFF0;
    // rom_array[26607] = 32'hFFFFFFF0;
    // rom_array[26608] = 32'hFFFFFFF0;
    // rom_array[26609] = 32'hFFFFFFF1;
    // rom_array[26610] = 32'hFFFFFFF1;
    // rom_array[26611] = 32'hFFFFFFF1;
    // rom_array[26612] = 32'hFFFFFFF1;
    // rom_array[26613] = 32'hFFFFFFF0;
    // rom_array[26614] = 32'hFFFFFFF0;
    // rom_array[26615] = 32'hFFFFFFF0;
    // rom_array[26616] = 32'hFFFFFFF0;
    // rom_array[26617] = 32'hFFFFFFF1;
    // rom_array[26618] = 32'hFFFFFFF1;
    // rom_array[26619] = 32'hFFFFFFF1;
    // rom_array[26620] = 32'hFFFFFFF1;
    // rom_array[26621] = 32'hFFFFFFF1;
    // rom_array[26622] = 32'hFFFFFFF1;
    // rom_array[26623] = 32'hFFFFFFF1;
    // rom_array[26624] = 32'hFFFFFFF1;
    // rom_array[26625] = 32'hFFFFFFF1;
    // rom_array[26626] = 32'hFFFFFFF1;
    // rom_array[26627] = 32'hFFFFFFF1;
    // rom_array[26628] = 32'hFFFFFFF1;
    // rom_array[26629] = 32'hFFFFFFF1;
    // rom_array[26630] = 32'hFFFFFFF1;
    // rom_array[26631] = 32'hFFFFFFF1;
    // rom_array[26632] = 32'hFFFFFFF1;
    // rom_array[26633] = 32'hFFFFFFF1;
    // rom_array[26634] = 32'hFFFFFFF1;
    // rom_array[26635] = 32'hFFFFFFF0;
    // rom_array[26636] = 32'hFFFFFFF0;
    // rom_array[26637] = 32'hFFFFFFF1;
    // rom_array[26638] = 32'hFFFFFFF1;
    // rom_array[26639] = 32'hFFFFFFF0;
    // rom_array[26640] = 32'hFFFFFFF0;
    // rom_array[26641] = 32'hFFFFFFF1;
    // rom_array[26642] = 32'hFFFFFFF1;
    // rom_array[26643] = 32'hFFFFFFF0;
    // rom_array[26644] = 32'hFFFFFFF0;
    // rom_array[26645] = 32'hFFFFFFF1;
    // rom_array[26646] = 32'hFFFFFFF1;
    // rom_array[26647] = 32'hFFFFFFF0;
    // rom_array[26648] = 32'hFFFFFFF0;
    // rom_array[26649] = 32'hFFFFFFF1;
    // rom_array[26650] = 32'hFFFFFFF1;
    // rom_array[26651] = 32'hFFFFFFF1;
    // rom_array[26652] = 32'hFFFFFFF1;
    // rom_array[26653] = 32'hFFFFFFF1;
    // rom_array[26654] = 32'hFFFFFFF1;
    // rom_array[26655] = 32'hFFFFFFF1;
    // rom_array[26656] = 32'hFFFFFFF1;
    // rom_array[26657] = 32'hFFFFFFF1;
    // rom_array[26658] = 32'hFFFFFFF1;
    // rom_array[26659] = 32'hFFFFFFF1;
    // rom_array[26660] = 32'hFFFFFFF1;
    // rom_array[26661] = 32'hFFFFFFF1;
    // rom_array[26662] = 32'hFFFFFFF1;
    // rom_array[26663] = 32'hFFFFFFF1;
    // rom_array[26664] = 32'hFFFFFFF1;
    // rom_array[26665] = 32'hFFFFFFF1;
    // rom_array[26666] = 32'hFFFFFFF1;
    // rom_array[26667] = 32'hFFFFFFF0;
    // rom_array[26668] = 32'hFFFFFFF0;
    // rom_array[26669] = 32'hFFFFFFF1;
    // rom_array[26670] = 32'hFFFFFFF1;
    // rom_array[26671] = 32'hFFFFFFF0;
    // rom_array[26672] = 32'hFFFFFFF0;
    // rom_array[26673] = 32'hFFFFFFF1;
    // rom_array[26674] = 32'hFFFFFFF1;
    // rom_array[26675] = 32'hFFFFFFF0;
    // rom_array[26676] = 32'hFFFFFFF0;
    // rom_array[26677] = 32'hFFFFFFF1;
    // rom_array[26678] = 32'hFFFFFFF1;
    // rom_array[26679] = 32'hFFFFFFF0;
    // rom_array[26680] = 32'hFFFFFFF0;
    // rom_array[26681] = 32'hFFFFFFF1;
    // rom_array[26682] = 32'hFFFFFFF1;
    // rom_array[26683] = 32'hFFFFFFF1;
    // rom_array[26684] = 32'hFFFFFFF1;
    // rom_array[26685] = 32'hFFFFFFF0;
    // rom_array[26686] = 32'hFFFFFFF0;
    // rom_array[26687] = 32'hFFFFFFF0;
    // rom_array[26688] = 32'hFFFFFFF0;
    // rom_array[26689] = 32'hFFFFFFF1;
    // rom_array[26690] = 32'hFFFFFFF1;
    // rom_array[26691] = 32'hFFFFFFF1;
    // rom_array[26692] = 32'hFFFFFFF1;
    // rom_array[26693] = 32'hFFFFFFF0;
    // rom_array[26694] = 32'hFFFFFFF0;
    // rom_array[26695] = 32'hFFFFFFF0;
    // rom_array[26696] = 32'hFFFFFFF0;
    // rom_array[26697] = 32'hFFFFFFF1;
    // rom_array[26698] = 32'hFFFFFFF1;
    // rom_array[26699] = 32'hFFFFFFF1;
    // rom_array[26700] = 32'hFFFFFFF1;
    // rom_array[26701] = 32'hFFFFFFF0;
    // rom_array[26702] = 32'hFFFFFFF0;
    // rom_array[26703] = 32'hFFFFFFF0;
    // rom_array[26704] = 32'hFFFFFFF0;
    // rom_array[26705] = 32'hFFFFFFF1;
    // rom_array[26706] = 32'hFFFFFFF1;
    // rom_array[26707] = 32'hFFFFFFF1;
    // rom_array[26708] = 32'hFFFFFFF1;
    // rom_array[26709] = 32'hFFFFFFF0;
    // rom_array[26710] = 32'hFFFFFFF0;
    // rom_array[26711] = 32'hFFFFFFF0;
    // rom_array[26712] = 32'hFFFFFFF0;
    // rom_array[26713] = 32'hFFFFFFF1;
    // rom_array[26714] = 32'hFFFFFFF1;
    // rom_array[26715] = 32'hFFFFFFF1;
    // rom_array[26716] = 32'hFFFFFFF1;
    // rom_array[26717] = 32'hFFFFFFF0;
    // rom_array[26718] = 32'hFFFFFFF0;
    // rom_array[26719] = 32'hFFFFFFF0;
    // rom_array[26720] = 32'hFFFFFFF0;
    // rom_array[26721] = 32'hFFFFFFF1;
    // rom_array[26722] = 32'hFFFFFFF1;
    // rom_array[26723] = 32'hFFFFFFF1;
    // rom_array[26724] = 32'hFFFFFFF1;
    // rom_array[26725] = 32'hFFFFFFF0;
    // rom_array[26726] = 32'hFFFFFFF0;
    // rom_array[26727] = 32'hFFFFFFF0;
    // rom_array[26728] = 32'hFFFFFFF0;
    // rom_array[26729] = 32'hFFFFFFF1;
    // rom_array[26730] = 32'hFFFFFFF1;
    // rom_array[26731] = 32'hFFFFFFF0;
    // rom_array[26732] = 32'hFFFFFFF0;
    // rom_array[26733] = 32'hFFFFFFF1;
    // rom_array[26734] = 32'hFFFFFFF1;
    // rom_array[26735] = 32'hFFFFFFF0;
    // rom_array[26736] = 32'hFFFFFFF0;
    // rom_array[26737] = 32'hFFFFFFF1;
    // rom_array[26738] = 32'hFFFFFFF1;
    // rom_array[26739] = 32'hFFFFFFF0;
    // rom_array[26740] = 32'hFFFFFFF0;
    // rom_array[26741] = 32'hFFFFFFF1;
    // rom_array[26742] = 32'hFFFFFFF1;
    // rom_array[26743] = 32'hFFFFFFF0;
    // rom_array[26744] = 32'hFFFFFFF0;
    // rom_array[26745] = 32'hFFFFFFF1;
    // rom_array[26746] = 32'hFFFFFFF1;
    // rom_array[26747] = 32'hFFFFFFF0;
    // rom_array[26748] = 32'hFFFFFFF0;
    // rom_array[26749] = 32'hFFFFFFF1;
    // rom_array[26750] = 32'hFFFFFFF1;
    // rom_array[26751] = 32'hFFFFFFF0;
    // rom_array[26752] = 32'hFFFFFFF0;
    // rom_array[26753] = 32'hFFFFFFF1;
    // rom_array[26754] = 32'hFFFFFFF1;
    // rom_array[26755] = 32'hFFFFFFF0;
    // rom_array[26756] = 32'hFFFFFFF0;
    // rom_array[26757] = 32'hFFFFFFF1;
    // rom_array[26758] = 32'hFFFFFFF1;
    // rom_array[26759] = 32'hFFFFFFF0;
    // rom_array[26760] = 32'hFFFFFFF0;
    // rom_array[26761] = 32'hFFFFFFF1;
    // rom_array[26762] = 32'hFFFFFFF1;
    // rom_array[26763] = 32'hFFFFFFF0;
    // rom_array[26764] = 32'hFFFFFFF0;
    // rom_array[26765] = 32'hFFFFFFF1;
    // rom_array[26766] = 32'hFFFFFFF1;
    // rom_array[26767] = 32'hFFFFFFF0;
    // rom_array[26768] = 32'hFFFFFFF0;
    // rom_array[26769] = 32'hFFFFFFF1;
    // rom_array[26770] = 32'hFFFFFFF1;
    // rom_array[26771] = 32'hFFFFFFF0;
    // rom_array[26772] = 32'hFFFFFFF0;
    // rom_array[26773] = 32'hFFFFFFF1;
    // rom_array[26774] = 32'hFFFFFFF1;
    // rom_array[26775] = 32'hFFFFFFF0;
    // rom_array[26776] = 32'hFFFFFFF0;
    // rom_array[26777] = 32'hFFFFFFF1;
    // rom_array[26778] = 32'hFFFFFFF1;
    // rom_array[26779] = 32'hFFFFFFF0;
    // rom_array[26780] = 32'hFFFFFFF0;
    // rom_array[26781] = 32'hFFFFFFF1;
    // rom_array[26782] = 32'hFFFFFFF1;
    // rom_array[26783] = 32'hFFFFFFF0;
    // rom_array[26784] = 32'hFFFFFFF0;
    // rom_array[26785] = 32'hFFFFFFF1;
    // rom_array[26786] = 32'hFFFFFFF1;
    // rom_array[26787] = 32'hFFFFFFF0;
    // rom_array[26788] = 32'hFFFFFFF0;
    // rom_array[26789] = 32'hFFFFFFF1;
    // rom_array[26790] = 32'hFFFFFFF1;
    // rom_array[26791] = 32'hFFFFFFF0;
    // rom_array[26792] = 32'hFFFFFFF0;
    // rom_array[26793] = 32'hFFFFFFF1;
    // rom_array[26794] = 32'hFFFFFFF1;
    // rom_array[26795] = 32'hFFFFFFF0;
    // rom_array[26796] = 32'hFFFFFFF0;
    // rom_array[26797] = 32'hFFFFFFF1;
    // rom_array[26798] = 32'hFFFFFFF1;
    // rom_array[26799] = 32'hFFFFFFF0;
    // rom_array[26800] = 32'hFFFFFFF0;
    // rom_array[26801] = 32'hFFFFFFF1;
    // rom_array[26802] = 32'hFFFFFFF1;
    // rom_array[26803] = 32'hFFFFFFF0;
    // rom_array[26804] = 32'hFFFFFFF0;
    // rom_array[26805] = 32'hFFFFFFF1;
    // rom_array[26806] = 32'hFFFFFFF1;
    // rom_array[26807] = 32'hFFFFFFF0;
    // rom_array[26808] = 32'hFFFFFFF0;
    // rom_array[26809] = 32'hFFFFFFF1;
    // rom_array[26810] = 32'hFFFFFFF1;
    // rom_array[26811] = 32'hFFFFFFF0;
    // rom_array[26812] = 32'hFFFFFFF0;
    // rom_array[26813] = 32'hFFFFFFF1;
    // rom_array[26814] = 32'hFFFFFFF1;
    // rom_array[26815] = 32'hFFFFFFF0;
    // rom_array[26816] = 32'hFFFFFFF0;
    // rom_array[26817] = 32'hFFFFFFF1;
    // rom_array[26818] = 32'hFFFFFFF1;
    // rom_array[26819] = 32'hFFFFFFF0;
    // rom_array[26820] = 32'hFFFFFFF0;
    // rom_array[26821] = 32'hFFFFFFF1;
    // rom_array[26822] = 32'hFFFFFFF1;
    // rom_array[26823] = 32'hFFFFFFF0;
    // rom_array[26824] = 32'hFFFFFFF0;
    // rom_array[26825] = 32'hFFFFFFF1;
    // rom_array[26826] = 32'hFFFFFFF1;
    // rom_array[26827] = 32'hFFFFFFF1;
    // rom_array[26828] = 32'hFFFFFFF1;
    // rom_array[26829] = 32'hFFFFFFF1;
    // rom_array[26830] = 32'hFFFFFFF1;
    // rom_array[26831] = 32'hFFFFFFF1;
    // rom_array[26832] = 32'hFFFFFFF1;
    // rom_array[26833] = 32'hFFFFFFF1;
    // rom_array[26834] = 32'hFFFFFFF1;
    // rom_array[26835] = 32'hFFFFFFF1;
    // rom_array[26836] = 32'hFFFFFFF1;
    // rom_array[26837] = 32'hFFFFFFF1;
    // rom_array[26838] = 32'hFFFFFFF1;
    // rom_array[26839] = 32'hFFFFFFF1;
    // rom_array[26840] = 32'hFFFFFFF1;
    // rom_array[26841] = 32'hFFFFFFF1;
    // rom_array[26842] = 32'hFFFFFFF1;
    // rom_array[26843] = 32'hFFFFFFF1;
    // rom_array[26844] = 32'hFFFFFFF1;
    // rom_array[26845] = 32'hFFFFFFF1;
    // rom_array[26846] = 32'hFFFFFFF1;
    // rom_array[26847] = 32'hFFFFFFF1;
    // rom_array[26848] = 32'hFFFFFFF1;
    // rom_array[26849] = 32'hFFFFFFF1;
    // rom_array[26850] = 32'hFFFFFFF1;
    // rom_array[26851] = 32'hFFFFFFF1;
    // rom_array[26852] = 32'hFFFFFFF1;
    // rom_array[26853] = 32'hFFFFFFF1;
    // rom_array[26854] = 32'hFFFFFFF1;
    // rom_array[26855] = 32'hFFFFFFF1;
    // rom_array[26856] = 32'hFFFFFFF1;
    // rom_array[26857] = 32'hFFFFFFF1;
    // rom_array[26858] = 32'hFFFFFFF1;
    // rom_array[26859] = 32'hFFFFFFF1;
    // rom_array[26860] = 32'hFFFFFFF1;
    // rom_array[26861] = 32'hFFFFFFF1;
    // rom_array[26862] = 32'hFFFFFFF1;
    // rom_array[26863] = 32'hFFFFFFF1;
    // rom_array[26864] = 32'hFFFFFFF1;
    // rom_array[26865] = 32'hFFFFFFF1;
    // rom_array[26866] = 32'hFFFFFFF1;
    // rom_array[26867] = 32'hFFFFFFF1;
    // rom_array[26868] = 32'hFFFFFFF1;
    // rom_array[26869] = 32'hFFFFFFF1;
    // rom_array[26870] = 32'hFFFFFFF1;
    // rom_array[26871] = 32'hFFFFFFF1;
    // rom_array[26872] = 32'hFFFFFFF1;
    // rom_array[26873] = 32'hFFFFFFF1;
    // rom_array[26874] = 32'hFFFFFFF1;
    // rom_array[26875] = 32'hFFFFFFF1;
    // rom_array[26876] = 32'hFFFFFFF1;
    // rom_array[26877] = 32'hFFFFFFF1;
    // rom_array[26878] = 32'hFFFFFFF1;
    // rom_array[26879] = 32'hFFFFFFF1;
    // rom_array[26880] = 32'hFFFFFFF1;
    // rom_array[26881] = 32'hFFFFFFF1;
    // rom_array[26882] = 32'hFFFFFFF1;
    // rom_array[26883] = 32'hFFFFFFF1;
    // rom_array[26884] = 32'hFFFFFFF1;
    // rom_array[26885] = 32'hFFFFFFF1;
    // rom_array[26886] = 32'hFFFFFFF1;
    // rom_array[26887] = 32'hFFFFFFF1;
    // rom_array[26888] = 32'hFFFFFFF1;
    // rom_array[26889] = 32'hFFFFFFF1;
    // rom_array[26890] = 32'hFFFFFFF1;
    // rom_array[26891] = 32'hFFFFFFF1;
    // rom_array[26892] = 32'hFFFFFFF1;
    // rom_array[26893] = 32'hFFFFFFF1;
    // rom_array[26894] = 32'hFFFFFFF1;
    // rom_array[26895] = 32'hFFFFFFF1;
    // rom_array[26896] = 32'hFFFFFFF1;
    // rom_array[26897] = 32'hFFFFFFF1;
    // rom_array[26898] = 32'hFFFFFFF1;
    // rom_array[26899] = 32'hFFFFFFF1;
    // rom_array[26900] = 32'hFFFFFFF1;
    // rom_array[26901] = 32'hFFFFFFF1;
    // rom_array[26902] = 32'hFFFFFFF1;
    // rom_array[26903] = 32'hFFFFFFF1;
    // rom_array[26904] = 32'hFFFFFFF1;
    // rom_array[26905] = 32'hFFFFFFF1;
    // rom_array[26906] = 32'hFFFFFFF1;
    // rom_array[26907] = 32'hFFFFFFF1;
    // rom_array[26908] = 32'hFFFFFFF1;
    // rom_array[26909] = 32'hFFFFFFF1;
    // rom_array[26910] = 32'hFFFFFFF1;
    // rom_array[26911] = 32'hFFFFFFF1;
    // rom_array[26912] = 32'hFFFFFFF1;
    // rom_array[26913] = 32'hFFFFFFF1;
    // rom_array[26914] = 32'hFFFFFFF1;
    // rom_array[26915] = 32'hFFFFFFF1;
    // rom_array[26916] = 32'hFFFFFFF1;
    // rom_array[26917] = 32'hFFFFFFF1;
    // rom_array[26918] = 32'hFFFFFFF1;
    // rom_array[26919] = 32'hFFFFFFF1;
    // rom_array[26920] = 32'hFFFFFFF1;
    // rom_array[26921] = 32'hFFFFFFF1;
    // rom_array[26922] = 32'hFFFFFFF1;
    // rom_array[26923] = 32'hFFFFFFF1;
    // rom_array[26924] = 32'hFFFFFFF1;
    // rom_array[26925] = 32'hFFFFFFF1;
    // rom_array[26926] = 32'hFFFFFFF1;
    // rom_array[26927] = 32'hFFFFFFF1;
    // rom_array[26928] = 32'hFFFFFFF1;
    // rom_array[26929] = 32'hFFFFFFF1;
    // rom_array[26930] = 32'hFFFFFFF1;
    // rom_array[26931] = 32'hFFFFFFF1;
    // rom_array[26932] = 32'hFFFFFFF1;
    // rom_array[26933] = 32'hFFFFFFF1;
    // rom_array[26934] = 32'hFFFFFFF1;
    // rom_array[26935] = 32'hFFFFFFF1;
    // rom_array[26936] = 32'hFFFFFFF1;
    // rom_array[26937] = 32'hFFFFFFF1;
    // rom_array[26938] = 32'hFFFFFFF1;
    // rom_array[26939] = 32'hFFFFFFF1;
    // rom_array[26940] = 32'hFFFFFFF1;
    // rom_array[26941] = 32'hFFFFFFF1;
    // rom_array[26942] = 32'hFFFFFFF1;
    // rom_array[26943] = 32'hFFFFFFF1;
    // rom_array[26944] = 32'hFFFFFFF1;
    // rom_array[26945] = 32'hFFFFFFF1;
    // rom_array[26946] = 32'hFFFFFFF1;
    // rom_array[26947] = 32'hFFFFFFF1;
    // rom_array[26948] = 32'hFFFFFFF1;
    // rom_array[26949] = 32'hFFFFFFF1;
    // rom_array[26950] = 32'hFFFFFFF1;
    // rom_array[26951] = 32'hFFFFFFF1;
    // rom_array[26952] = 32'hFFFFFFF1;
    // rom_array[26953] = 32'hFFFFFFF1;
    // rom_array[26954] = 32'hFFFFFFF1;
    // rom_array[26955] = 32'hFFFFFFF1;
    // rom_array[26956] = 32'hFFFFFFF1;
    // rom_array[26957] = 32'hFFFFFFF1;
    // rom_array[26958] = 32'hFFFFFFF1;
    // rom_array[26959] = 32'hFFFFFFF1;
    // rom_array[26960] = 32'hFFFFFFF1;
    // rom_array[26961] = 32'hFFFFFFF1;
    // rom_array[26962] = 32'hFFFFFFF1;
    // rom_array[26963] = 32'hFFFFFFF1;
    // rom_array[26964] = 32'hFFFFFFF1;
    // rom_array[26965] = 32'hFFFFFFF1;
    // rom_array[26966] = 32'hFFFFFFF1;
    // rom_array[26967] = 32'hFFFFFFF1;
    // rom_array[26968] = 32'hFFFFFFF1;
    // rom_array[26969] = 32'hFFFFFFF1;
    // rom_array[26970] = 32'hFFFFFFF1;
    // rom_array[26971] = 32'hFFFFFFF1;
    // rom_array[26972] = 32'hFFFFFFF1;
    // rom_array[26973] = 32'hFFFFFFF1;
    // rom_array[26974] = 32'hFFFFFFF1;
    // rom_array[26975] = 32'hFFFFFFF1;
    // rom_array[26976] = 32'hFFFFFFF1;
    // rom_array[26977] = 32'hFFFFFFF1;
    // rom_array[26978] = 32'hFFFFFFF1;
    // rom_array[26979] = 32'hFFFFFFF1;
    // rom_array[26980] = 32'hFFFFFFF1;
    // rom_array[26981] = 32'hFFFFFFF1;
    // rom_array[26982] = 32'hFFFFFFF1;
    // rom_array[26983] = 32'hFFFFFFF1;
    // rom_array[26984] = 32'hFFFFFFF1;
    // rom_array[26985] = 32'hFFFFFFF1;
    // rom_array[26986] = 32'hFFFFFFF1;
    // rom_array[26987] = 32'hFFFFFFF1;
    // rom_array[26988] = 32'hFFFFFFF1;
    // rom_array[26989] = 32'hFFFFFFF1;
    // rom_array[26990] = 32'hFFFFFFF1;
    // rom_array[26991] = 32'hFFFFFFF1;
    // rom_array[26992] = 32'hFFFFFFF1;
    // rom_array[26993] = 32'hFFFFFFF1;
    // rom_array[26994] = 32'hFFFFFFF1;
    // rom_array[26995] = 32'hFFFFFFF1;
    // rom_array[26996] = 32'hFFFFFFF1;
    // rom_array[26997] = 32'hFFFFFFF1;
    // rom_array[26998] = 32'hFFFFFFF1;
    // rom_array[26999] = 32'hFFFFFFF1;
    // rom_array[27000] = 32'hFFFFFFF1;
    // rom_array[27001] = 32'hFFFFFFF1;
    // rom_array[27002] = 32'hFFFFFFF1;
    // rom_array[27003] = 32'hFFFFFFF1;
    // rom_array[27004] = 32'hFFFFFFF1;
    // rom_array[27005] = 32'hFFFFFFF1;
    // rom_array[27006] = 32'hFFFFFFF1;
    // rom_array[27007] = 32'hFFFFFFF1;
    // rom_array[27008] = 32'hFFFFFFF1;
    // rom_array[27009] = 32'hFFFFFFF1;
    // rom_array[27010] = 32'hFFFFFFF1;
    // rom_array[27011] = 32'hFFFFFFF1;
    // rom_array[27012] = 32'hFFFFFFF1;
    // rom_array[27013] = 32'hFFFFFFF1;
    // rom_array[27014] = 32'hFFFFFFF1;
    // rom_array[27015] = 32'hFFFFFFF1;
    // rom_array[27016] = 32'hFFFFFFF1;
    // rom_array[27017] = 32'hFFFFFFF1;
    // rom_array[27018] = 32'hFFFFFFF1;
    // rom_array[27019] = 32'hFFFFFFF1;
    // rom_array[27020] = 32'hFFFFFFF1;
    // rom_array[27021] = 32'hFFFFFFF1;
    // rom_array[27022] = 32'hFFFFFFF1;
    // rom_array[27023] = 32'hFFFFFFF1;
    // rom_array[27024] = 32'hFFFFFFF1;
    // rom_array[27025] = 32'hFFFFFFF1;
    // rom_array[27026] = 32'hFFFFFFF1;
    // rom_array[27027] = 32'hFFFFFFF1;
    // rom_array[27028] = 32'hFFFFFFF1;
    // rom_array[27029] = 32'hFFFFFFF1;
    // rom_array[27030] = 32'hFFFFFFF1;
    // rom_array[27031] = 32'hFFFFFFF1;
    // rom_array[27032] = 32'hFFFFFFF1;
    // rom_array[27033] = 32'hFFFFFFF1;
    // rom_array[27034] = 32'hFFFFFFF1;
    // rom_array[27035] = 32'hFFFFFFF1;
    // rom_array[27036] = 32'hFFFFFFF1;
    // rom_array[27037] = 32'hFFFFFFF1;
    // rom_array[27038] = 32'hFFFFFFF1;
    // rom_array[27039] = 32'hFFFFFFF1;
    // rom_array[27040] = 32'hFFFFFFF1;
    // rom_array[27041] = 32'hFFFFFFF1;
    // rom_array[27042] = 32'hFFFFFFF1;
    // rom_array[27043] = 32'hFFFFFFF1;
    // rom_array[27044] = 32'hFFFFFFF1;
    // rom_array[27045] = 32'hFFFFFFF1;
    // rom_array[27046] = 32'hFFFFFFF1;
    // rom_array[27047] = 32'hFFFFFFF1;
    // rom_array[27048] = 32'hFFFFFFF1;
    // rom_array[27049] = 32'hFFFFFFF1;
    // rom_array[27050] = 32'hFFFFFFF1;
    // rom_array[27051] = 32'hFFFFFFF1;
    // rom_array[27052] = 32'hFFFFFFF1;
    // rom_array[27053] = 32'hFFFFFFF1;
    // rom_array[27054] = 32'hFFFFFFF1;
    // rom_array[27055] = 32'hFFFFFFF1;
    // rom_array[27056] = 32'hFFFFFFF1;
    // rom_array[27057] = 32'hFFFFFFF1;
    // rom_array[27058] = 32'hFFFFFFF1;
    // rom_array[27059] = 32'hFFFFFFF1;
    // rom_array[27060] = 32'hFFFFFFF1;
    // rom_array[27061] = 32'hFFFFFFF1;
    // rom_array[27062] = 32'hFFFFFFF1;
    // rom_array[27063] = 32'hFFFFFFF1;
    // rom_array[27064] = 32'hFFFFFFF1;
    // rom_array[27065] = 32'hFFFFFFF1;
    // rom_array[27066] = 32'hFFFFFFF1;
    // rom_array[27067] = 32'hFFFFFFF1;
    // rom_array[27068] = 32'hFFFFFFF1;
    // rom_array[27069] = 32'hFFFFFFF1;
    // rom_array[27070] = 32'hFFFFFFF1;
    // rom_array[27071] = 32'hFFFFFFF1;
    // rom_array[27072] = 32'hFFFFFFF1;
    // rom_array[27073] = 32'hFFFFFFF1;
    // rom_array[27074] = 32'hFFFFFFF1;
    // rom_array[27075] = 32'hFFFFFFF1;
    // rom_array[27076] = 32'hFFFFFFF1;
    // rom_array[27077] = 32'hFFFFFFF1;
    // rom_array[27078] = 32'hFFFFFFF1;
    // rom_array[27079] = 32'hFFFFFFF1;
    // rom_array[27080] = 32'hFFFFFFF1;
    // rom_array[27081] = 32'hFFFFFFF1;
    // rom_array[27082] = 32'hFFFFFFF1;
    // rom_array[27083] = 32'hFFFFFFF1;
    // rom_array[27084] = 32'hFFFFFFF1;
    // rom_array[27085] = 32'hFFFFFFF1;
    // rom_array[27086] = 32'hFFFFFFF1;
    // rom_array[27087] = 32'hFFFFFFF1;
    // rom_array[27088] = 32'hFFFFFFF1;
    // rom_array[27089] = 32'hFFFFFFF1;
    // rom_array[27090] = 32'hFFFFFFF1;
    // rom_array[27091] = 32'hFFFFFFF1;
    // rom_array[27092] = 32'hFFFFFFF1;
    // rom_array[27093] = 32'hFFFFFFF1;
    // rom_array[27094] = 32'hFFFFFFF1;
    // rom_array[27095] = 32'hFFFFFFF1;
    // rom_array[27096] = 32'hFFFFFFF1;
    // rom_array[27097] = 32'hFFFFFFF1;
    // rom_array[27098] = 32'hFFFFFFF1;
    // rom_array[27099] = 32'hFFFFFFF1;
    // rom_array[27100] = 32'hFFFFFFF1;
    // rom_array[27101] = 32'hFFFFFFF1;
    // rom_array[27102] = 32'hFFFFFFF1;
    // rom_array[27103] = 32'hFFFFFFF1;
    // rom_array[27104] = 32'hFFFFFFF1;
    // rom_array[27105] = 32'hFFFFFFF1;
    // rom_array[27106] = 32'hFFFFFFF1;
    // rom_array[27107] = 32'hFFFFFFF1;
    // rom_array[27108] = 32'hFFFFFFF1;
    // rom_array[27109] = 32'hFFFFFFF1;
    // rom_array[27110] = 32'hFFFFFFF1;
    // rom_array[27111] = 32'hFFFFFFF1;
    // rom_array[27112] = 32'hFFFFFFF1;
    // rom_array[27113] = 32'hFFFFFFF1;
    // rom_array[27114] = 32'hFFFFFFF1;
    // rom_array[27115] = 32'hFFFFFFF1;
    // rom_array[27116] = 32'hFFFFFFF1;
    // rom_array[27117] = 32'hFFFFFFF1;
    // rom_array[27118] = 32'hFFFFFFF1;
    // rom_array[27119] = 32'hFFFFFFF1;
    // rom_array[27120] = 32'hFFFFFFF1;
    // rom_array[27121] = 32'hFFFFFFF1;
    // rom_array[27122] = 32'hFFFFFFF1;
    // rom_array[27123] = 32'hFFFFFFF1;
    // rom_array[27124] = 32'hFFFFFFF1;
    // rom_array[27125] = 32'hFFFFFFF1;
    // rom_array[27126] = 32'hFFFFFFF1;
    // rom_array[27127] = 32'hFFFFFFF1;
    // rom_array[27128] = 32'hFFFFFFF1;
    // rom_array[27129] = 32'hFFFFFFF1;
    // rom_array[27130] = 32'hFFFFFFF1;
    // rom_array[27131] = 32'hFFFFFFF0;
    // rom_array[27132] = 32'hFFFFFFF0;
    // rom_array[27133] = 32'hFFFFFFF1;
    // rom_array[27134] = 32'hFFFFFFF1;
    // rom_array[27135] = 32'hFFFFFFF0;
    // rom_array[27136] = 32'hFFFFFFF0;
    // rom_array[27137] = 32'hFFFFFFF1;
    // rom_array[27138] = 32'hFFFFFFF1;
    // rom_array[27139] = 32'hFFFFFFF0;
    // rom_array[27140] = 32'hFFFFFFF0;
    // rom_array[27141] = 32'hFFFFFFF1;
    // rom_array[27142] = 32'hFFFFFFF1;
    // rom_array[27143] = 32'hFFFFFFF0;
    // rom_array[27144] = 32'hFFFFFFF0;
    // rom_array[27145] = 32'hFFFFFFF1;
    // rom_array[27146] = 32'hFFFFFFF1;
    // rom_array[27147] = 32'hFFFFFFF0;
    // rom_array[27148] = 32'hFFFFFFF0;
    // rom_array[27149] = 32'hFFFFFFF1;
    // rom_array[27150] = 32'hFFFFFFF1;
    // rom_array[27151] = 32'hFFFFFFF0;
    // rom_array[27152] = 32'hFFFFFFF0;
    // rom_array[27153] = 32'hFFFFFFF1;
    // rom_array[27154] = 32'hFFFFFFF1;
    // rom_array[27155] = 32'hFFFFFFF0;
    // rom_array[27156] = 32'hFFFFFFF0;
    // rom_array[27157] = 32'hFFFFFFF1;
    // rom_array[27158] = 32'hFFFFFFF1;
    // rom_array[27159] = 32'hFFFFFFF0;
    // rom_array[27160] = 32'hFFFFFFF0;
    // rom_array[27161] = 32'hFFFFFFF1;
    // rom_array[27162] = 32'hFFFFFFF1;
    // rom_array[27163] = 32'hFFFFFFF1;
    // rom_array[27164] = 32'hFFFFFFF1;
    // rom_array[27165] = 32'hFFFFFFF1;
    // rom_array[27166] = 32'hFFFFFFF1;
    // rom_array[27167] = 32'hFFFFFFF1;
    // rom_array[27168] = 32'hFFFFFFF1;
    // rom_array[27169] = 32'hFFFFFFF1;
    // rom_array[27170] = 32'hFFFFFFF1;
    // rom_array[27171] = 32'hFFFFFFF1;
    // rom_array[27172] = 32'hFFFFFFF1;
    // rom_array[27173] = 32'hFFFFFFF1;
    // rom_array[27174] = 32'hFFFFFFF1;
    // rom_array[27175] = 32'hFFFFFFF1;
    // rom_array[27176] = 32'hFFFFFFF1;
    // rom_array[27177] = 32'hFFFFFFF1;
    // rom_array[27178] = 32'hFFFFFFF1;
    // rom_array[27179] = 32'hFFFFFFF1;
    // rom_array[27180] = 32'hFFFFFFF1;
    // rom_array[27181] = 32'hFFFFFFF1;
    // rom_array[27182] = 32'hFFFFFFF1;
    // rom_array[27183] = 32'hFFFFFFF1;
    // rom_array[27184] = 32'hFFFFFFF1;
    // rom_array[27185] = 32'hFFFFFFF1;
    // rom_array[27186] = 32'hFFFFFFF1;
    // rom_array[27187] = 32'hFFFFFFF1;
    // rom_array[27188] = 32'hFFFFFFF1;
    // rom_array[27189] = 32'hFFFFFFF1;
    // rom_array[27190] = 32'hFFFFFFF1;
    // rom_array[27191] = 32'hFFFFFFF1;
    // rom_array[27192] = 32'hFFFFFFF1;
    // rom_array[27193] = 32'hFFFFFFF1;
    // rom_array[27194] = 32'hFFFFFFF1;
    // rom_array[27195] = 32'hFFFFFFF1;
    // rom_array[27196] = 32'hFFFFFFF1;
    // rom_array[27197] = 32'hFFFFFFF1;
    // rom_array[27198] = 32'hFFFFFFF1;
    // rom_array[27199] = 32'hFFFFFFF1;
    // rom_array[27200] = 32'hFFFFFFF1;
    // rom_array[27201] = 32'hFFFFFFF1;
    // rom_array[27202] = 32'hFFFFFFF1;
    // rom_array[27203] = 32'hFFFFFFF1;
    // rom_array[27204] = 32'hFFFFFFF1;
    // rom_array[27205] = 32'hFFFFFFF1;
    // rom_array[27206] = 32'hFFFFFFF1;
    // rom_array[27207] = 32'hFFFFFFF1;
    // rom_array[27208] = 32'hFFFFFFF1;
    // rom_array[27209] = 32'hFFFFFFF1;
    // rom_array[27210] = 32'hFFFFFFF1;
    // rom_array[27211] = 32'hFFFFFFF0;
    // rom_array[27212] = 32'hFFFFFFF0;
    // rom_array[27213] = 32'hFFFFFFF1;
    // rom_array[27214] = 32'hFFFFFFF1;
    // rom_array[27215] = 32'hFFFFFFF0;
    // rom_array[27216] = 32'hFFFFFFF0;
    // rom_array[27217] = 32'hFFFFFFF1;
    // rom_array[27218] = 32'hFFFFFFF1;
    // rom_array[27219] = 32'hFFFFFFF0;
    // rom_array[27220] = 32'hFFFFFFF0;
    // rom_array[27221] = 32'hFFFFFFF1;
    // rom_array[27222] = 32'hFFFFFFF1;
    // rom_array[27223] = 32'hFFFFFFF0;
    // rom_array[27224] = 32'hFFFFFFF0;
    // rom_array[27225] = 32'hFFFFFFF1;
    // rom_array[27226] = 32'hFFFFFFF1;
    // rom_array[27227] = 32'hFFFFFFF0;
    // rom_array[27228] = 32'hFFFFFFF0;
    // rom_array[27229] = 32'hFFFFFFF1;
    // rom_array[27230] = 32'hFFFFFFF1;
    // rom_array[27231] = 32'hFFFFFFF0;
    // rom_array[27232] = 32'hFFFFFFF0;
    // rom_array[27233] = 32'hFFFFFFF1;
    // rom_array[27234] = 32'hFFFFFFF1;
    // rom_array[27235] = 32'hFFFFFFF0;
    // rom_array[27236] = 32'hFFFFFFF0;
    // rom_array[27237] = 32'hFFFFFFF1;
    // rom_array[27238] = 32'hFFFFFFF1;
    // rom_array[27239] = 32'hFFFFFFF0;
    // rom_array[27240] = 32'hFFFFFFF0;
    // rom_array[27241] = 32'hFFFFFFF1;
    // rom_array[27242] = 32'hFFFFFFF1;
    // rom_array[27243] = 32'hFFFFFFF0;
    // rom_array[27244] = 32'hFFFFFFF0;
    // rom_array[27245] = 32'hFFFFFFF1;
    // rom_array[27246] = 32'hFFFFFFF1;
    // rom_array[27247] = 32'hFFFFFFF0;
    // rom_array[27248] = 32'hFFFFFFF0;
    // rom_array[27249] = 32'hFFFFFFF1;
    // rom_array[27250] = 32'hFFFFFFF1;
    // rom_array[27251] = 32'hFFFFFFF0;
    // rom_array[27252] = 32'hFFFFFFF0;
    // rom_array[27253] = 32'hFFFFFFF1;
    // rom_array[27254] = 32'hFFFFFFF1;
    // rom_array[27255] = 32'hFFFFFFF0;
    // rom_array[27256] = 32'hFFFFFFF0;
    // rom_array[27257] = 32'hFFFFFFF1;
    // rom_array[27258] = 32'hFFFFFFF1;
    // rom_array[27259] = 32'hFFFFFFF0;
    // rom_array[27260] = 32'hFFFFFFF0;
    // rom_array[27261] = 32'hFFFFFFF1;
    // rom_array[27262] = 32'hFFFFFFF1;
    // rom_array[27263] = 32'hFFFFFFF0;
    // rom_array[27264] = 32'hFFFFFFF0;
    // rom_array[27265] = 32'hFFFFFFF1;
    // rom_array[27266] = 32'hFFFFFFF1;
    // rom_array[27267] = 32'hFFFFFFF0;
    // rom_array[27268] = 32'hFFFFFFF0;
    // rom_array[27269] = 32'hFFFFFFF1;
    // rom_array[27270] = 32'hFFFFFFF1;
    // rom_array[27271] = 32'hFFFFFFF0;
    // rom_array[27272] = 32'hFFFFFFF0;
    // rom_array[27273] = 32'hFFFFFFF1;
    // rom_array[27274] = 32'hFFFFFFF1;
    // rom_array[27275] = 32'hFFFFFFF0;
    // rom_array[27276] = 32'hFFFFFFF0;
    // rom_array[27277] = 32'hFFFFFFF1;
    // rom_array[27278] = 32'hFFFFFFF1;
    // rom_array[27279] = 32'hFFFFFFF0;
    // rom_array[27280] = 32'hFFFFFFF0;
    // rom_array[27281] = 32'hFFFFFFF1;
    // rom_array[27282] = 32'hFFFFFFF1;
    // rom_array[27283] = 32'hFFFFFFF0;
    // rom_array[27284] = 32'hFFFFFFF0;
    // rom_array[27285] = 32'hFFFFFFF1;
    // rom_array[27286] = 32'hFFFFFFF1;
    // rom_array[27287] = 32'hFFFFFFF0;
    // rom_array[27288] = 32'hFFFFFFF0;
    // rom_array[27289] = 32'hFFFFFFF1;
    // rom_array[27290] = 32'hFFFFFFF1;
    // rom_array[27291] = 32'hFFFFFFF0;
    // rom_array[27292] = 32'hFFFFFFF0;
    // rom_array[27293] = 32'hFFFFFFF1;
    // rom_array[27294] = 32'hFFFFFFF1;
    // rom_array[27295] = 32'hFFFFFFF0;
    // rom_array[27296] = 32'hFFFFFFF0;
    // rom_array[27297] = 32'hFFFFFFF1;
    // rom_array[27298] = 32'hFFFFFFF1;
    // rom_array[27299] = 32'hFFFFFFF0;
    // rom_array[27300] = 32'hFFFFFFF0;
    // rom_array[27301] = 32'hFFFFFFF1;
    // rom_array[27302] = 32'hFFFFFFF1;
    // rom_array[27303] = 32'hFFFFFFF0;
    // rom_array[27304] = 32'hFFFFFFF0;
    // rom_array[27305] = 32'hFFFFFFF0;
    // rom_array[27306] = 32'hFFFFFFF0;
    // rom_array[27307] = 32'hFFFFFFF0;
    // rom_array[27308] = 32'hFFFFFFF0;
    // rom_array[27309] = 32'hFFFFFFF1;
    // rom_array[27310] = 32'hFFFFFFF1;
    // rom_array[27311] = 32'hFFFFFFF1;
    // rom_array[27312] = 32'hFFFFFFF1;
    // rom_array[27313] = 32'hFFFFFFF0;
    // rom_array[27314] = 32'hFFFFFFF0;
    // rom_array[27315] = 32'hFFFFFFF0;
    // rom_array[27316] = 32'hFFFFFFF0;
    // rom_array[27317] = 32'hFFFFFFF1;
    // rom_array[27318] = 32'hFFFFFFF1;
    // rom_array[27319] = 32'hFFFFFFF1;
    // rom_array[27320] = 32'hFFFFFFF1;
    // rom_array[27321] = 32'hFFFFFFF0;
    // rom_array[27322] = 32'hFFFFFFF0;
    // rom_array[27323] = 32'hFFFFFFF0;
    // rom_array[27324] = 32'hFFFFFFF0;
    // rom_array[27325] = 32'hFFFFFFF1;
    // rom_array[27326] = 32'hFFFFFFF1;
    // rom_array[27327] = 32'hFFFFFFF1;
    // rom_array[27328] = 32'hFFFFFFF1;
    // rom_array[27329] = 32'hFFFFFFF0;
    // rom_array[27330] = 32'hFFFFFFF0;
    // rom_array[27331] = 32'hFFFFFFF0;
    // rom_array[27332] = 32'hFFFFFFF0;
    // rom_array[27333] = 32'hFFFFFFF1;
    // rom_array[27334] = 32'hFFFFFFF1;
    // rom_array[27335] = 32'hFFFFFFF1;
    // rom_array[27336] = 32'hFFFFFFF1;
    // rom_array[27337] = 32'hFFFFFFF0;
    // rom_array[27338] = 32'hFFFFFFF0;
    // rom_array[27339] = 32'hFFFFFFF0;
    // rom_array[27340] = 32'hFFFFFFF0;
    // rom_array[27341] = 32'hFFFFFFF1;
    // rom_array[27342] = 32'hFFFFFFF1;
    // rom_array[27343] = 32'hFFFFFFF1;
    // rom_array[27344] = 32'hFFFFFFF1;
    // rom_array[27345] = 32'hFFFFFFF0;
    // rom_array[27346] = 32'hFFFFFFF0;
    // rom_array[27347] = 32'hFFFFFFF0;
    // rom_array[27348] = 32'hFFFFFFF0;
    // rom_array[27349] = 32'hFFFFFFF1;
    // rom_array[27350] = 32'hFFFFFFF1;
    // rom_array[27351] = 32'hFFFFFFF1;
    // rom_array[27352] = 32'hFFFFFFF1;
    // rom_array[27353] = 32'hFFFFFFF0;
    // rom_array[27354] = 32'hFFFFFFF0;
    // rom_array[27355] = 32'hFFFFFFF0;
    // rom_array[27356] = 32'hFFFFFFF0;
    // rom_array[27357] = 32'hFFFFFFF1;
    // rom_array[27358] = 32'hFFFFFFF1;
    // rom_array[27359] = 32'hFFFFFFF1;
    // rom_array[27360] = 32'hFFFFFFF1;
    // rom_array[27361] = 32'hFFFFFFF0;
    // rom_array[27362] = 32'hFFFFFFF0;
    // rom_array[27363] = 32'hFFFFFFF0;
    // rom_array[27364] = 32'hFFFFFFF0;
    // rom_array[27365] = 32'hFFFFFFF1;
    // rom_array[27366] = 32'hFFFFFFF1;
    // rom_array[27367] = 32'hFFFFFFF1;
    // rom_array[27368] = 32'hFFFFFFF1;
    // rom_array[27369] = 32'hFFFFFFF1;
    // rom_array[27370] = 32'hFFFFFFF1;
    // rom_array[27371] = 32'hFFFFFFF1;
    // rom_array[27372] = 32'hFFFFFFF1;
    // rom_array[27373] = 32'hFFFFFFF1;
    // rom_array[27374] = 32'hFFFFFFF1;
    // rom_array[27375] = 32'hFFFFFFF1;
    // rom_array[27376] = 32'hFFFFFFF1;
    // rom_array[27377] = 32'hFFFFFFF1;
    // rom_array[27378] = 32'hFFFFFFF1;
    // rom_array[27379] = 32'hFFFFFFF1;
    // rom_array[27380] = 32'hFFFFFFF1;
    // rom_array[27381] = 32'hFFFFFFF1;
    // rom_array[27382] = 32'hFFFFFFF1;
    // rom_array[27383] = 32'hFFFFFFF1;
    // rom_array[27384] = 32'hFFFFFFF1;
    // rom_array[27385] = 32'hFFFFFFF1;
    // rom_array[27386] = 32'hFFFFFFF1;
    // rom_array[27387] = 32'hFFFFFFF1;
    // rom_array[27388] = 32'hFFFFFFF1;
    // rom_array[27389] = 32'hFFFFFFF1;
    // rom_array[27390] = 32'hFFFFFFF1;
    // rom_array[27391] = 32'hFFFFFFF1;
    // rom_array[27392] = 32'hFFFFFFF1;
    // rom_array[27393] = 32'hFFFFFFF1;
    // rom_array[27394] = 32'hFFFFFFF1;
    // rom_array[27395] = 32'hFFFFFFF1;
    // rom_array[27396] = 32'hFFFFFFF1;
    // rom_array[27397] = 32'hFFFFFFF1;
    // rom_array[27398] = 32'hFFFFFFF1;
    // rom_array[27399] = 32'hFFFFFFF1;
    // rom_array[27400] = 32'hFFFFFFF1;
    // rom_array[27401] = 32'hFFFFFFF1;
    // rom_array[27402] = 32'hFFFFFFF1;
    // rom_array[27403] = 32'hFFFFFFF1;
    // rom_array[27404] = 32'hFFFFFFF1;
    // rom_array[27405] = 32'hFFFFFFF1;
    // rom_array[27406] = 32'hFFFFFFF1;
    // rom_array[27407] = 32'hFFFFFFF1;
    // rom_array[27408] = 32'hFFFFFFF1;
    // rom_array[27409] = 32'hFFFFFFF1;
    // rom_array[27410] = 32'hFFFFFFF1;
    // rom_array[27411] = 32'hFFFFFFF1;
    // rom_array[27412] = 32'hFFFFFFF1;
    // rom_array[27413] = 32'hFFFFFFF1;
    // rom_array[27414] = 32'hFFFFFFF1;
    // rom_array[27415] = 32'hFFFFFFF1;
    // rom_array[27416] = 32'hFFFFFFF1;
    // rom_array[27417] = 32'hFFFFFFF1;
    // rom_array[27418] = 32'hFFFFFFF1;
    // rom_array[27419] = 32'hFFFFFFF1;
    // rom_array[27420] = 32'hFFFFFFF1;
    // rom_array[27421] = 32'hFFFFFFF1;
    // rom_array[27422] = 32'hFFFFFFF1;
    // rom_array[27423] = 32'hFFFFFFF1;
    // rom_array[27424] = 32'hFFFFFFF1;
    // rom_array[27425] = 32'hFFFFFFF1;
    // rom_array[27426] = 32'hFFFFFFF1;
    // rom_array[27427] = 32'hFFFFFFF1;
    // rom_array[27428] = 32'hFFFFFFF1;
    // rom_array[27429] = 32'hFFFFFFF1;
    // rom_array[27430] = 32'hFFFFFFF1;
    // rom_array[27431] = 32'hFFFFFFF1;
    // rom_array[27432] = 32'hFFFFFFF1;
    // rom_array[27433] = 32'hFFFFFFF0;
    // rom_array[27434] = 32'hFFFFFFF0;
    // rom_array[27435] = 32'hFFFFFFF0;
    // rom_array[27436] = 32'hFFFFFFF0;
    // rom_array[27437] = 32'hFFFFFFF1;
    // rom_array[27438] = 32'hFFFFFFF1;
    // rom_array[27439] = 32'hFFFFFFF1;
    // rom_array[27440] = 32'hFFFFFFF1;
    // rom_array[27441] = 32'hFFFFFFF0;
    // rom_array[27442] = 32'hFFFFFFF0;
    // rom_array[27443] = 32'hFFFFFFF0;
    // rom_array[27444] = 32'hFFFFFFF0;
    // rom_array[27445] = 32'hFFFFFFF1;
    // rom_array[27446] = 32'hFFFFFFF1;
    // rom_array[27447] = 32'hFFFFFFF1;
    // rom_array[27448] = 32'hFFFFFFF1;
    // rom_array[27449] = 32'hFFFFFFF0;
    // rom_array[27450] = 32'hFFFFFFF0;
    // rom_array[27451] = 32'hFFFFFFF0;
    // rom_array[27452] = 32'hFFFFFFF0;
    // rom_array[27453] = 32'hFFFFFFF1;
    // rom_array[27454] = 32'hFFFFFFF1;
    // rom_array[27455] = 32'hFFFFFFF1;
    // rom_array[27456] = 32'hFFFFFFF1;
    // rom_array[27457] = 32'hFFFFFFF0;
    // rom_array[27458] = 32'hFFFFFFF0;
    // rom_array[27459] = 32'hFFFFFFF0;
    // rom_array[27460] = 32'hFFFFFFF0;
    // rom_array[27461] = 32'hFFFFFFF1;
    // rom_array[27462] = 32'hFFFFFFF1;
    // rom_array[27463] = 32'hFFFFFFF1;
    // rom_array[27464] = 32'hFFFFFFF1;
    // rom_array[27465] = 32'hFFFFFFF0;
    // rom_array[27466] = 32'hFFFFFFF0;
    // rom_array[27467] = 32'hFFFFFFF0;
    // rom_array[27468] = 32'hFFFFFFF0;
    // rom_array[27469] = 32'hFFFFFFF1;
    // rom_array[27470] = 32'hFFFFFFF1;
    // rom_array[27471] = 32'hFFFFFFF1;
    // rom_array[27472] = 32'hFFFFFFF1;
    // rom_array[27473] = 32'hFFFFFFF0;
    // rom_array[27474] = 32'hFFFFFFF0;
    // rom_array[27475] = 32'hFFFFFFF0;
    // rom_array[27476] = 32'hFFFFFFF0;
    // rom_array[27477] = 32'hFFFFFFF1;
    // rom_array[27478] = 32'hFFFFFFF1;
    // rom_array[27479] = 32'hFFFFFFF1;
    // rom_array[27480] = 32'hFFFFFFF1;
    // rom_array[27481] = 32'hFFFFFFF0;
    // rom_array[27482] = 32'hFFFFFFF0;
    // rom_array[27483] = 32'hFFFFFFF0;
    // rom_array[27484] = 32'hFFFFFFF0;
    // rom_array[27485] = 32'hFFFFFFF1;
    // rom_array[27486] = 32'hFFFFFFF1;
    // rom_array[27487] = 32'hFFFFFFF1;
    // rom_array[27488] = 32'hFFFFFFF1;
    // rom_array[27489] = 32'hFFFFFFF0;
    // rom_array[27490] = 32'hFFFFFFF0;
    // rom_array[27491] = 32'hFFFFFFF0;
    // rom_array[27492] = 32'hFFFFFFF0;
    // rom_array[27493] = 32'hFFFFFFF1;
    // rom_array[27494] = 32'hFFFFFFF1;
    // rom_array[27495] = 32'hFFFFFFF1;
    // rom_array[27496] = 32'hFFFFFFF1;
    // rom_array[27497] = 32'hFFFFFFF1;
    // rom_array[27498] = 32'hFFFFFFF1;
    // rom_array[27499] = 32'hFFFFFFF1;
    // rom_array[27500] = 32'hFFFFFFF1;
    // rom_array[27501] = 32'hFFFFFFF1;
    // rom_array[27502] = 32'hFFFFFFF1;
    // rom_array[27503] = 32'hFFFFFFF1;
    // rom_array[27504] = 32'hFFFFFFF1;
    // rom_array[27505] = 32'hFFFFFFF1;
    // rom_array[27506] = 32'hFFFFFFF1;
    // rom_array[27507] = 32'hFFFFFFF1;
    // rom_array[27508] = 32'hFFFFFFF1;
    // rom_array[27509] = 32'hFFFFFFF1;
    // rom_array[27510] = 32'hFFFFFFF1;
    // rom_array[27511] = 32'hFFFFFFF1;
    // rom_array[27512] = 32'hFFFFFFF1;
    // rom_array[27513] = 32'hFFFFFFF1;
    // rom_array[27514] = 32'hFFFFFFF1;
    // rom_array[27515] = 32'hFFFFFFF1;
    // rom_array[27516] = 32'hFFFFFFF1;
    // rom_array[27517] = 32'hFFFFFFF1;
    // rom_array[27518] = 32'hFFFFFFF1;
    // rom_array[27519] = 32'hFFFFFFF1;
    // rom_array[27520] = 32'hFFFFFFF1;
    // rom_array[27521] = 32'hFFFFFFF1;
    // rom_array[27522] = 32'hFFFFFFF1;
    // rom_array[27523] = 32'hFFFFFFF1;
    // rom_array[27524] = 32'hFFFFFFF1;
    // rom_array[27525] = 32'hFFFFFFF1;
    // rom_array[27526] = 32'hFFFFFFF1;
    // rom_array[27527] = 32'hFFFFFFF1;
    // rom_array[27528] = 32'hFFFFFFF1;
    // rom_array[27529] = 32'hFFFFFFF1;
    // rom_array[27530] = 32'hFFFFFFF1;
    // rom_array[27531] = 32'hFFFFFFF1;
    // rom_array[27532] = 32'hFFFFFFF1;
    // rom_array[27533] = 32'hFFFFFFF1;
    // rom_array[27534] = 32'hFFFFFFF1;
    // rom_array[27535] = 32'hFFFFFFF1;
    // rom_array[27536] = 32'hFFFFFFF1;
    // rom_array[27537] = 32'hFFFFFFF1;
    // rom_array[27538] = 32'hFFFFFFF1;
    // rom_array[27539] = 32'hFFFFFFF1;
    // rom_array[27540] = 32'hFFFFFFF1;
    // rom_array[27541] = 32'hFFFFFFF1;
    // rom_array[27542] = 32'hFFFFFFF1;
    // rom_array[27543] = 32'hFFFFFFF1;
    // rom_array[27544] = 32'hFFFFFFF1;
    // rom_array[27545] = 32'hFFFFFFF1;
    // rom_array[27546] = 32'hFFFFFFF1;
    // rom_array[27547] = 32'hFFFFFFF1;
    // rom_array[27548] = 32'hFFFFFFF1;
    // rom_array[27549] = 32'hFFFFFFF1;
    // rom_array[27550] = 32'hFFFFFFF1;
    // rom_array[27551] = 32'hFFFFFFF1;
    // rom_array[27552] = 32'hFFFFFFF1;
    // rom_array[27553] = 32'hFFFFFFF1;
    // rom_array[27554] = 32'hFFFFFFF1;
    // rom_array[27555] = 32'hFFFFFFF1;
    // rom_array[27556] = 32'hFFFFFFF1;
    // rom_array[27557] = 32'hFFFFFFF1;
    // rom_array[27558] = 32'hFFFFFFF1;
    // rom_array[27559] = 32'hFFFFFFF1;
    // rom_array[27560] = 32'hFFFFFFF1;
    // rom_array[27561] = 32'hFFFFFFF1;
    // rom_array[27562] = 32'hFFFFFFF1;
    // rom_array[27563] = 32'hFFFFFFF1;
    // rom_array[27564] = 32'hFFFFFFF1;
    // rom_array[27565] = 32'hFFFFFFF0;
    // rom_array[27566] = 32'hFFFFFFF0;
    // rom_array[27567] = 32'hFFFFFFF0;
    // rom_array[27568] = 32'hFFFFFFF0;
    // rom_array[27569] = 32'hFFFFFFF1;
    // rom_array[27570] = 32'hFFFFFFF1;
    // rom_array[27571] = 32'hFFFFFFF1;
    // rom_array[27572] = 32'hFFFFFFF1;
    // rom_array[27573] = 32'hFFFFFFF0;
    // rom_array[27574] = 32'hFFFFFFF0;
    // rom_array[27575] = 32'hFFFFFFF0;
    // rom_array[27576] = 32'hFFFFFFF0;
    // rom_array[27577] = 32'hFFFFFFF1;
    // rom_array[27578] = 32'hFFFFFFF1;
    // rom_array[27579] = 32'hFFFFFFF1;
    // rom_array[27580] = 32'hFFFFFFF1;
    // rom_array[27581] = 32'hFFFFFFF0;
    // rom_array[27582] = 32'hFFFFFFF0;
    // rom_array[27583] = 32'hFFFFFFF0;
    // rom_array[27584] = 32'hFFFFFFF0;
    // rom_array[27585] = 32'hFFFFFFF1;
    // rom_array[27586] = 32'hFFFFFFF1;
    // rom_array[27587] = 32'hFFFFFFF1;
    // rom_array[27588] = 32'hFFFFFFF1;
    // rom_array[27589] = 32'hFFFFFFF0;
    // rom_array[27590] = 32'hFFFFFFF0;
    // rom_array[27591] = 32'hFFFFFFF0;
    // rom_array[27592] = 32'hFFFFFFF0;
    // rom_array[27593] = 32'hFFFFFFF1;
    // rom_array[27594] = 32'hFFFFFFF1;
    // rom_array[27595] = 32'hFFFFFFF1;
    // rom_array[27596] = 32'hFFFFFFF1;
    // rom_array[27597] = 32'hFFFFFFF0;
    // rom_array[27598] = 32'hFFFFFFF0;
    // rom_array[27599] = 32'hFFFFFFF0;
    // rom_array[27600] = 32'hFFFFFFF0;
    // rom_array[27601] = 32'hFFFFFFF1;
    // rom_array[27602] = 32'hFFFFFFF1;
    // rom_array[27603] = 32'hFFFFFFF1;
    // rom_array[27604] = 32'hFFFFFFF1;
    // rom_array[27605] = 32'hFFFFFFF0;
    // rom_array[27606] = 32'hFFFFFFF0;
    // rom_array[27607] = 32'hFFFFFFF0;
    // rom_array[27608] = 32'hFFFFFFF0;
    // rom_array[27609] = 32'hFFFFFFF1;
    // rom_array[27610] = 32'hFFFFFFF1;
    // rom_array[27611] = 32'hFFFFFFF1;
    // rom_array[27612] = 32'hFFFFFFF1;
    // rom_array[27613] = 32'hFFFFFFF0;
    // rom_array[27614] = 32'hFFFFFFF0;
    // rom_array[27615] = 32'hFFFFFFF0;
    // rom_array[27616] = 32'hFFFFFFF0;
    // rom_array[27617] = 32'hFFFFFFF1;
    // rom_array[27618] = 32'hFFFFFFF1;
    // rom_array[27619] = 32'hFFFFFFF1;
    // rom_array[27620] = 32'hFFFFFFF1;
    // rom_array[27621] = 32'hFFFFFFF0;
    // rom_array[27622] = 32'hFFFFFFF0;
    // rom_array[27623] = 32'hFFFFFFF0;
    // rom_array[27624] = 32'hFFFFFFF0;
    // rom_array[27625] = 32'hFFFFFFF1;
    // rom_array[27626] = 32'hFFFFFFF1;
    // rom_array[27627] = 32'hFFFFFFF1;
    // rom_array[27628] = 32'hFFFFFFF1;
    // rom_array[27629] = 32'hFFFFFFF0;
    // rom_array[27630] = 32'hFFFFFFF0;
    // rom_array[27631] = 32'hFFFFFFF0;
    // rom_array[27632] = 32'hFFFFFFF0;
    // rom_array[27633] = 32'hFFFFFFF1;
    // rom_array[27634] = 32'hFFFFFFF1;
    // rom_array[27635] = 32'hFFFFFFF1;
    // rom_array[27636] = 32'hFFFFFFF1;
    // rom_array[27637] = 32'hFFFFFFF0;
    // rom_array[27638] = 32'hFFFFFFF0;
    // rom_array[27639] = 32'hFFFFFFF0;
    // rom_array[27640] = 32'hFFFFFFF0;
    // rom_array[27641] = 32'hFFFFFFF1;
    // rom_array[27642] = 32'hFFFFFFF1;
    // rom_array[27643] = 32'hFFFFFFF1;
    // rom_array[27644] = 32'hFFFFFFF1;
    // rom_array[27645] = 32'hFFFFFFF0;
    // rom_array[27646] = 32'hFFFFFFF0;
    // rom_array[27647] = 32'hFFFFFFF0;
    // rom_array[27648] = 32'hFFFFFFF0;
    // rom_array[27649] = 32'hFFFFFFF1;
    // rom_array[27650] = 32'hFFFFFFF1;
    // rom_array[27651] = 32'hFFFFFFF1;
    // rom_array[27652] = 32'hFFFFFFF1;
    // rom_array[27653] = 32'hFFFFFFF0;
    // rom_array[27654] = 32'hFFFFFFF0;
    // rom_array[27655] = 32'hFFFFFFF0;
    // rom_array[27656] = 32'hFFFFFFF0;
    // rom_array[27657] = 32'hFFFFFFF1;
    // rom_array[27658] = 32'hFFFFFFF1;
    // rom_array[27659] = 32'hFFFFFFF1;
    // rom_array[27660] = 32'hFFFFFFF1;
    // rom_array[27661] = 32'hFFFFFFF0;
    // rom_array[27662] = 32'hFFFFFFF0;
    // rom_array[27663] = 32'hFFFFFFF0;
    // rom_array[27664] = 32'hFFFFFFF0;
    // rom_array[27665] = 32'hFFFFFFF1;
    // rom_array[27666] = 32'hFFFFFFF1;
    // rom_array[27667] = 32'hFFFFFFF1;
    // rom_array[27668] = 32'hFFFFFFF1;
    // rom_array[27669] = 32'hFFFFFFF0;
    // rom_array[27670] = 32'hFFFFFFF0;
    // rom_array[27671] = 32'hFFFFFFF0;
    // rom_array[27672] = 32'hFFFFFFF0;
    // rom_array[27673] = 32'hFFFFFFF1;
    // rom_array[27674] = 32'hFFFFFFF1;
    // rom_array[27675] = 32'hFFFFFFF1;
    // rom_array[27676] = 32'hFFFFFFF1;
    // rom_array[27677] = 32'hFFFFFFF0;
    // rom_array[27678] = 32'hFFFFFFF0;
    // rom_array[27679] = 32'hFFFFFFF0;
    // rom_array[27680] = 32'hFFFFFFF0;
    // rom_array[27681] = 32'hFFFFFFF1;
    // rom_array[27682] = 32'hFFFFFFF1;
    // rom_array[27683] = 32'hFFFFFFF1;
    // rom_array[27684] = 32'hFFFFFFF1;
    // rom_array[27685] = 32'hFFFFFFF0;
    // rom_array[27686] = 32'hFFFFFFF0;
    // rom_array[27687] = 32'hFFFFFFF0;
    // rom_array[27688] = 32'hFFFFFFF0;
    // rom_array[27689] = 32'hFFFFFFF0;
    // rom_array[27690] = 32'hFFFFFFF0;
    // rom_array[27691] = 32'hFFFFFFF0;
    // rom_array[27692] = 32'hFFFFFFF0;
    // rom_array[27693] = 32'hFFFFFFF1;
    // rom_array[27694] = 32'hFFFFFFF1;
    // rom_array[27695] = 32'hFFFFFFF1;
    // rom_array[27696] = 32'hFFFFFFF1;
    // rom_array[27697] = 32'hFFFFFFF0;
    // rom_array[27698] = 32'hFFFFFFF0;
    // rom_array[27699] = 32'hFFFFFFF0;
    // rom_array[27700] = 32'hFFFFFFF0;
    // rom_array[27701] = 32'hFFFFFFF1;
    // rom_array[27702] = 32'hFFFFFFF1;
    // rom_array[27703] = 32'hFFFFFFF1;
    // rom_array[27704] = 32'hFFFFFFF1;
    // rom_array[27705] = 32'hFFFFFFF0;
    // rom_array[27706] = 32'hFFFFFFF0;
    // rom_array[27707] = 32'hFFFFFFF0;
    // rom_array[27708] = 32'hFFFFFFF0;
    // rom_array[27709] = 32'hFFFFFFF1;
    // rom_array[27710] = 32'hFFFFFFF1;
    // rom_array[27711] = 32'hFFFFFFF1;
    // rom_array[27712] = 32'hFFFFFFF1;
    // rom_array[27713] = 32'hFFFFFFF0;
    // rom_array[27714] = 32'hFFFFFFF0;
    // rom_array[27715] = 32'hFFFFFFF0;
    // rom_array[27716] = 32'hFFFFFFF0;
    // rom_array[27717] = 32'hFFFFFFF1;
    // rom_array[27718] = 32'hFFFFFFF1;
    // rom_array[27719] = 32'hFFFFFFF1;
    // rom_array[27720] = 32'hFFFFFFF1;
    // rom_array[27721] = 32'hFFFFFFF0;
    // rom_array[27722] = 32'hFFFFFFF0;
    // rom_array[27723] = 32'hFFFFFFF0;
    // rom_array[27724] = 32'hFFFFFFF0;
    // rom_array[27725] = 32'hFFFFFFF1;
    // rom_array[27726] = 32'hFFFFFFF1;
    // rom_array[27727] = 32'hFFFFFFF1;
    // rom_array[27728] = 32'hFFFFFFF1;
    // rom_array[27729] = 32'hFFFFFFF0;
    // rom_array[27730] = 32'hFFFFFFF0;
    // rom_array[27731] = 32'hFFFFFFF0;
    // rom_array[27732] = 32'hFFFFFFF0;
    // rom_array[27733] = 32'hFFFFFFF1;
    // rom_array[27734] = 32'hFFFFFFF1;
    // rom_array[27735] = 32'hFFFFFFF1;
    // rom_array[27736] = 32'hFFFFFFF1;
    // rom_array[27737] = 32'hFFFFFFF1;
    // rom_array[27738] = 32'hFFFFFFF1;
    // rom_array[27739] = 32'hFFFFFFF0;
    // rom_array[27740] = 32'hFFFFFFF0;
    // rom_array[27741] = 32'hFFFFFFF1;
    // rom_array[27742] = 32'hFFFFFFF1;
    // rom_array[27743] = 32'hFFFFFFF0;
    // rom_array[27744] = 32'hFFFFFFF0;
    // rom_array[27745] = 32'hFFFFFFF1;
    // rom_array[27746] = 32'hFFFFFFF1;
    // rom_array[27747] = 32'hFFFFFFF0;
    // rom_array[27748] = 32'hFFFFFFF0;
    // rom_array[27749] = 32'hFFFFFFF1;
    // rom_array[27750] = 32'hFFFFFFF1;
    // rom_array[27751] = 32'hFFFFFFF0;
    // rom_array[27752] = 32'hFFFFFFF0;
    // rom_array[27753] = 32'hFFFFFFF1;
    // rom_array[27754] = 32'hFFFFFFF1;
    // rom_array[27755] = 32'hFFFFFFF1;
    // rom_array[27756] = 32'hFFFFFFF1;
    // rom_array[27757] = 32'hFFFFFFF1;
    // rom_array[27758] = 32'hFFFFFFF1;
    // rom_array[27759] = 32'hFFFFFFF1;
    // rom_array[27760] = 32'hFFFFFFF1;
    // rom_array[27761] = 32'hFFFFFFF1;
    // rom_array[27762] = 32'hFFFFFFF1;
    // rom_array[27763] = 32'hFFFFFFF1;
    // rom_array[27764] = 32'hFFFFFFF1;
    // rom_array[27765] = 32'hFFFFFFF1;
    // rom_array[27766] = 32'hFFFFFFF1;
    // rom_array[27767] = 32'hFFFFFFF1;
    // rom_array[27768] = 32'hFFFFFFF1;
    // rom_array[27769] = 32'hFFFFFFF1;
    // rom_array[27770] = 32'hFFFFFFF1;
    // rom_array[27771] = 32'hFFFFFFF0;
    // rom_array[27772] = 32'hFFFFFFF0;
    // rom_array[27773] = 32'hFFFFFFF1;
    // rom_array[27774] = 32'hFFFFFFF1;
    // rom_array[27775] = 32'hFFFFFFF0;
    // rom_array[27776] = 32'hFFFFFFF0;
    // rom_array[27777] = 32'hFFFFFFF1;
    // rom_array[27778] = 32'hFFFFFFF1;
    // rom_array[27779] = 32'hFFFFFFF0;
    // rom_array[27780] = 32'hFFFFFFF0;
    // rom_array[27781] = 32'hFFFFFFF1;
    // rom_array[27782] = 32'hFFFFFFF1;
    // rom_array[27783] = 32'hFFFFFFF0;
    // rom_array[27784] = 32'hFFFFFFF0;
    // rom_array[27785] = 32'hFFFFFFF1;
    // rom_array[27786] = 32'hFFFFFFF1;
    // rom_array[27787] = 32'hFFFFFFF1;
    // rom_array[27788] = 32'hFFFFFFF1;
    // rom_array[27789] = 32'hFFFFFFF1;
    // rom_array[27790] = 32'hFFFFFFF1;
    // rom_array[27791] = 32'hFFFFFFF1;
    // rom_array[27792] = 32'hFFFFFFF1;
    // rom_array[27793] = 32'hFFFFFFF1;
    // rom_array[27794] = 32'hFFFFFFF1;
    // rom_array[27795] = 32'hFFFFFFF1;
    // rom_array[27796] = 32'hFFFFFFF1;
    // rom_array[27797] = 32'hFFFFFFF1;
    // rom_array[27798] = 32'hFFFFFFF1;
    // rom_array[27799] = 32'hFFFFFFF1;
    // rom_array[27800] = 32'hFFFFFFF1;
    // rom_array[27801] = 32'hFFFFFFF1;
    // rom_array[27802] = 32'hFFFFFFF1;
    // rom_array[27803] = 32'hFFFFFFF1;
    // rom_array[27804] = 32'hFFFFFFF1;
    // rom_array[27805] = 32'hFFFFFFF1;
    // rom_array[27806] = 32'hFFFFFFF1;
    // rom_array[27807] = 32'hFFFFFFF1;
    // rom_array[27808] = 32'hFFFFFFF1;
    // rom_array[27809] = 32'hFFFFFFF1;
    // rom_array[27810] = 32'hFFFFFFF1;
    // rom_array[27811] = 32'hFFFFFFF1;
    // rom_array[27812] = 32'hFFFFFFF1;
    // rom_array[27813] = 32'hFFFFFFF1;
    // rom_array[27814] = 32'hFFFFFFF1;
    // rom_array[27815] = 32'hFFFFFFF1;
    // rom_array[27816] = 32'hFFFFFFF1;
    // rom_array[27817] = 32'hFFFFFFF1;
    // rom_array[27818] = 32'hFFFFFFF1;
    // rom_array[27819] = 32'hFFFFFFF1;
    // rom_array[27820] = 32'hFFFFFFF1;
    // rom_array[27821] = 32'hFFFFFFF1;
    // rom_array[27822] = 32'hFFFFFFF1;
    // rom_array[27823] = 32'hFFFFFFF1;
    // rom_array[27824] = 32'hFFFFFFF1;
    // rom_array[27825] = 32'hFFFFFFF1;
    // rom_array[27826] = 32'hFFFFFFF1;
    // rom_array[27827] = 32'hFFFFFFF1;
    // rom_array[27828] = 32'hFFFFFFF1;
    // rom_array[27829] = 32'hFFFFFFF1;
    // rom_array[27830] = 32'hFFFFFFF1;
    // rom_array[27831] = 32'hFFFFFFF1;
    // rom_array[27832] = 32'hFFFFFFF1;
    // rom_array[27833] = 32'hFFFFFFF1;
    // rom_array[27834] = 32'hFFFFFFF1;
    // rom_array[27835] = 32'hFFFFFFF0;
    // rom_array[27836] = 32'hFFFFFFF0;
    // rom_array[27837] = 32'hFFFFFFF1;
    // rom_array[27838] = 32'hFFFFFFF1;
    // rom_array[27839] = 32'hFFFFFFF0;
    // rom_array[27840] = 32'hFFFFFFF0;
    // rom_array[27841] = 32'hFFFFFFF1;
    // rom_array[27842] = 32'hFFFFFFF1;
    // rom_array[27843] = 32'hFFFFFFF0;
    // rom_array[27844] = 32'hFFFFFFF0;
    // rom_array[27845] = 32'hFFFFFFF1;
    // rom_array[27846] = 32'hFFFFFFF1;
    // rom_array[27847] = 32'hFFFFFFF0;
    // rom_array[27848] = 32'hFFFFFFF0;
    // rom_array[27849] = 32'hFFFFFFF1;
    // rom_array[27850] = 32'hFFFFFFF1;
    // rom_array[27851] = 32'hFFFFFFF1;
    // rom_array[27852] = 32'hFFFFFFF1;
    // rom_array[27853] = 32'hFFFFFFF1;
    // rom_array[27854] = 32'hFFFFFFF1;
    // rom_array[27855] = 32'hFFFFFFF1;
    // rom_array[27856] = 32'hFFFFFFF1;
    // rom_array[27857] = 32'hFFFFFFF1;
    // rom_array[27858] = 32'hFFFFFFF1;
    // rom_array[27859] = 32'hFFFFFFF1;
    // rom_array[27860] = 32'hFFFFFFF1;
    // rom_array[27861] = 32'hFFFFFFF1;
    // rom_array[27862] = 32'hFFFFFFF1;
    // rom_array[27863] = 32'hFFFFFFF1;
    // rom_array[27864] = 32'hFFFFFFF1;
    // rom_array[27865] = 32'hFFFFFFF1;
    // rom_array[27866] = 32'hFFFFFFF1;
    // rom_array[27867] = 32'hFFFFFFF0;
    // rom_array[27868] = 32'hFFFFFFF0;
    // rom_array[27869] = 32'hFFFFFFF1;
    // rom_array[27870] = 32'hFFFFFFF1;
    // rom_array[27871] = 32'hFFFFFFF0;
    // rom_array[27872] = 32'hFFFFFFF0;
    // rom_array[27873] = 32'hFFFFFFF1;
    // rom_array[27874] = 32'hFFFFFFF1;
    // rom_array[27875] = 32'hFFFFFFF0;
    // rom_array[27876] = 32'hFFFFFFF0;
    // rom_array[27877] = 32'hFFFFFFF1;
    // rom_array[27878] = 32'hFFFFFFF1;
    // rom_array[27879] = 32'hFFFFFFF0;
    // rom_array[27880] = 32'hFFFFFFF0;
    // rom_array[27881] = 32'hFFFFFFF1;
    // rom_array[27882] = 32'hFFFFFFF1;
    // rom_array[27883] = 32'hFFFFFFF1;
    // rom_array[27884] = 32'hFFFFFFF1;
    // rom_array[27885] = 32'hFFFFFFF0;
    // rom_array[27886] = 32'hFFFFFFF0;
    // rom_array[27887] = 32'hFFFFFFF0;
    // rom_array[27888] = 32'hFFFFFFF0;
    // rom_array[27889] = 32'hFFFFFFF1;
    // rom_array[27890] = 32'hFFFFFFF1;
    // rom_array[27891] = 32'hFFFFFFF1;
    // rom_array[27892] = 32'hFFFFFFF1;
    // rom_array[27893] = 32'hFFFFFFF0;
    // rom_array[27894] = 32'hFFFFFFF0;
    // rom_array[27895] = 32'hFFFFFFF0;
    // rom_array[27896] = 32'hFFFFFFF0;
    // rom_array[27897] = 32'hFFFFFFF1;
    // rom_array[27898] = 32'hFFFFFFF1;
    // rom_array[27899] = 32'hFFFFFFF1;
    // rom_array[27900] = 32'hFFFFFFF1;
    // rom_array[27901] = 32'hFFFFFFF0;
    // rom_array[27902] = 32'hFFFFFFF0;
    // rom_array[27903] = 32'hFFFFFFF0;
    // rom_array[27904] = 32'hFFFFFFF0;
    // rom_array[27905] = 32'hFFFFFFF1;
    // rom_array[27906] = 32'hFFFFFFF1;
    // rom_array[27907] = 32'hFFFFFFF1;
    // rom_array[27908] = 32'hFFFFFFF1;
    // rom_array[27909] = 32'hFFFFFFF0;
    // rom_array[27910] = 32'hFFFFFFF0;
    // rom_array[27911] = 32'hFFFFFFF0;
    // rom_array[27912] = 32'hFFFFFFF0;
    // rom_array[27913] = 32'hFFFFFFF1;
    // rom_array[27914] = 32'hFFFFFFF1;
    // rom_array[27915] = 32'hFFFFFFF1;
    // rom_array[27916] = 32'hFFFFFFF1;
    // rom_array[27917] = 32'hFFFFFFF0;
    // rom_array[27918] = 32'hFFFFFFF0;
    // rom_array[27919] = 32'hFFFFFFF0;
    // rom_array[27920] = 32'hFFFFFFF0;
    // rom_array[27921] = 32'hFFFFFFF1;
    // rom_array[27922] = 32'hFFFFFFF1;
    // rom_array[27923] = 32'hFFFFFFF1;
    // rom_array[27924] = 32'hFFFFFFF1;
    // rom_array[27925] = 32'hFFFFFFF0;
    // rom_array[27926] = 32'hFFFFFFF0;
    // rom_array[27927] = 32'hFFFFFFF0;
    // rom_array[27928] = 32'hFFFFFFF0;
    // rom_array[27929] = 32'hFFFFFFF0;
    // rom_array[27930] = 32'hFFFFFFF0;
    // rom_array[27931] = 32'hFFFFFFF0;
    // rom_array[27932] = 32'hFFFFFFF0;
    // rom_array[27933] = 32'hFFFFFFF1;
    // rom_array[27934] = 32'hFFFFFFF1;
    // rom_array[27935] = 32'hFFFFFFF1;
    // rom_array[27936] = 32'hFFFFFFF1;
    // rom_array[27937] = 32'hFFFFFFF0;
    // rom_array[27938] = 32'hFFFFFFF0;
    // rom_array[27939] = 32'hFFFFFFF0;
    // rom_array[27940] = 32'hFFFFFFF0;
    // rom_array[27941] = 32'hFFFFFFF1;
    // rom_array[27942] = 32'hFFFFFFF1;
    // rom_array[27943] = 32'hFFFFFFF1;
    // rom_array[27944] = 32'hFFFFFFF1;
    // rom_array[27945] = 32'hFFFFFFF0;
    // rom_array[27946] = 32'hFFFFFFF0;
    // rom_array[27947] = 32'hFFFFFFF0;
    // rom_array[27948] = 32'hFFFFFFF0;
    // rom_array[27949] = 32'hFFFFFFF1;
    // rom_array[27950] = 32'hFFFFFFF1;
    // rom_array[27951] = 32'hFFFFFFF1;
    // rom_array[27952] = 32'hFFFFFFF1;
    // rom_array[27953] = 32'hFFFFFFF0;
    // rom_array[27954] = 32'hFFFFFFF0;
    // rom_array[27955] = 32'hFFFFFFF0;
    // rom_array[27956] = 32'hFFFFFFF0;
    // rom_array[27957] = 32'hFFFFFFF1;
    // rom_array[27958] = 32'hFFFFFFF1;
    // rom_array[27959] = 32'hFFFFFFF1;
    // rom_array[27960] = 32'hFFFFFFF1;
    // rom_array[27961] = 32'hFFFFFFF0;
    // rom_array[27962] = 32'hFFFFFFF0;
    // rom_array[27963] = 32'hFFFFFFF0;
    // rom_array[27964] = 32'hFFFFFFF0;
    // rom_array[27965] = 32'hFFFFFFF1;
    // rom_array[27966] = 32'hFFFFFFF1;
    // rom_array[27967] = 32'hFFFFFFF1;
    // rom_array[27968] = 32'hFFFFFFF1;
    // rom_array[27969] = 32'hFFFFFFF0;
    // rom_array[27970] = 32'hFFFFFFF0;
    // rom_array[27971] = 32'hFFFFFFF0;
    // rom_array[27972] = 32'hFFFFFFF0;
    // rom_array[27973] = 32'hFFFFFFF1;
    // rom_array[27974] = 32'hFFFFFFF1;
    // rom_array[27975] = 32'hFFFFFFF1;
    // rom_array[27976] = 32'hFFFFFFF1;
    // rom_array[27977] = 32'hFFFFFFF0;
    // rom_array[27978] = 32'hFFFFFFF0;
    // rom_array[27979] = 32'hFFFFFFF0;
    // rom_array[27980] = 32'hFFFFFFF0;
    // rom_array[27981] = 32'hFFFFFFF1;
    // rom_array[27982] = 32'hFFFFFFF1;
    // rom_array[27983] = 32'hFFFFFFF1;
    // rom_array[27984] = 32'hFFFFFFF1;
    // rom_array[27985] = 32'hFFFFFFF0;
    // rom_array[27986] = 32'hFFFFFFF0;
    // rom_array[27987] = 32'hFFFFFFF0;
    // rom_array[27988] = 32'hFFFFFFF0;
    // rom_array[27989] = 32'hFFFFFFF1;
    // rom_array[27990] = 32'hFFFFFFF1;
    // rom_array[27991] = 32'hFFFFFFF1;
    // rom_array[27992] = 32'hFFFFFFF1;
    // rom_array[27993] = 32'hFFFFFFF0;
    // rom_array[27994] = 32'hFFFFFFF0;
    // rom_array[27995] = 32'hFFFFFFF0;
    // rom_array[27996] = 32'hFFFFFFF0;
    // rom_array[27997] = 32'hFFFFFFF1;
    // rom_array[27998] = 32'hFFFFFFF1;
    // rom_array[27999] = 32'hFFFFFFF1;
    // rom_array[28000] = 32'hFFFFFFF1;
    // rom_array[28001] = 32'hFFFFFFF0;
    // rom_array[28002] = 32'hFFFFFFF0;
    // rom_array[28003] = 32'hFFFFFFF0;
    // rom_array[28004] = 32'hFFFFFFF0;
    // rom_array[28005] = 32'hFFFFFFF1;
    // rom_array[28006] = 32'hFFFFFFF1;
    // rom_array[28007] = 32'hFFFFFFF1;
    // rom_array[28008] = 32'hFFFFFFF1;
    // rom_array[28009] = 32'hFFFFFFF0;
    // rom_array[28010] = 32'hFFFFFFF0;
    // rom_array[28011] = 32'hFFFFFFF0;
    // rom_array[28012] = 32'hFFFFFFF0;
    // rom_array[28013] = 32'hFFFFFFF1;
    // rom_array[28014] = 32'hFFFFFFF1;
    // rom_array[28015] = 32'hFFFFFFF1;
    // rom_array[28016] = 32'hFFFFFFF1;
    // rom_array[28017] = 32'hFFFFFFF0;
    // rom_array[28018] = 32'hFFFFFFF0;
    // rom_array[28019] = 32'hFFFFFFF0;
    // rom_array[28020] = 32'hFFFFFFF0;
    // rom_array[28021] = 32'hFFFFFFF1;
    // rom_array[28022] = 32'hFFFFFFF1;
    // rom_array[28023] = 32'hFFFFFFF1;
    // rom_array[28024] = 32'hFFFFFFF1;
    // rom_array[28025] = 32'hFFFFFFF0;
    // rom_array[28026] = 32'hFFFFFFF0;
    // rom_array[28027] = 32'hFFFFFFF0;
    // rom_array[28028] = 32'hFFFFFFF0;
    // rom_array[28029] = 32'hFFFFFFF1;
    // rom_array[28030] = 32'hFFFFFFF1;
    // rom_array[28031] = 32'hFFFFFFF1;
    // rom_array[28032] = 32'hFFFFFFF1;
    // rom_array[28033] = 32'hFFFFFFF0;
    // rom_array[28034] = 32'hFFFFFFF0;
    // rom_array[28035] = 32'hFFFFFFF0;
    // rom_array[28036] = 32'hFFFFFFF0;
    // rom_array[28037] = 32'hFFFFFFF1;
    // rom_array[28038] = 32'hFFFFFFF1;
    // rom_array[28039] = 32'hFFFFFFF1;
    // rom_array[28040] = 32'hFFFFFFF1;
    // rom_array[28041] = 32'hFFFFFFF0;
    // rom_array[28042] = 32'hFFFFFFF0;
    // rom_array[28043] = 32'hFFFFFFF0;
    // rom_array[28044] = 32'hFFFFFFF0;
    // rom_array[28045] = 32'hFFFFFFF1;
    // rom_array[28046] = 32'hFFFFFFF1;
    // rom_array[28047] = 32'hFFFFFFF1;
    // rom_array[28048] = 32'hFFFFFFF1;
    // rom_array[28049] = 32'hFFFFFFF0;
    // rom_array[28050] = 32'hFFFFFFF0;
    // rom_array[28051] = 32'hFFFFFFF0;
    // rom_array[28052] = 32'hFFFFFFF0;
    // rom_array[28053] = 32'hFFFFFFF1;
    // rom_array[28054] = 32'hFFFFFFF1;
    // rom_array[28055] = 32'hFFFFFFF1;
    // rom_array[28056] = 32'hFFFFFFF1;
    // rom_array[28057] = 32'hFFFFFFF1;
    // rom_array[28058] = 32'hFFFFFFF1;
    // rom_array[28059] = 32'hFFFFFFF1;
    // rom_array[28060] = 32'hFFFFFFF1;
    // rom_array[28061] = 32'hFFFFFFF1;
    // rom_array[28062] = 32'hFFFFFFF1;
    // rom_array[28063] = 32'hFFFFFFF1;
    // rom_array[28064] = 32'hFFFFFFF1;
    // rom_array[28065] = 32'hFFFFFFF1;
    // rom_array[28066] = 32'hFFFFFFF1;
    // rom_array[28067] = 32'hFFFFFFF1;
    // rom_array[28068] = 32'hFFFFFFF1;
    // rom_array[28069] = 32'hFFFFFFF1;
    // rom_array[28070] = 32'hFFFFFFF1;
    // rom_array[28071] = 32'hFFFFFFF1;
    // rom_array[28072] = 32'hFFFFFFF1;
    // rom_array[28073] = 32'hFFFFFFF1;
    // rom_array[28074] = 32'hFFFFFFF1;
    // rom_array[28075] = 32'hFFFFFFF1;
    // rom_array[28076] = 32'hFFFFFFF1;
    // rom_array[28077] = 32'hFFFFFFF0;
    // rom_array[28078] = 32'hFFFFFFF0;
    // rom_array[28079] = 32'hFFFFFFF0;
    // rom_array[28080] = 32'hFFFFFFF0;
    // rom_array[28081] = 32'hFFFFFFF1;
    // rom_array[28082] = 32'hFFFFFFF1;
    // rom_array[28083] = 32'hFFFFFFF1;
    // rom_array[28084] = 32'hFFFFFFF1;
    // rom_array[28085] = 32'hFFFFFFF0;
    // rom_array[28086] = 32'hFFFFFFF0;
    // rom_array[28087] = 32'hFFFFFFF0;
    // rom_array[28088] = 32'hFFFFFFF0;
    // rom_array[28089] = 32'hFFFFFFF1;
    // rom_array[28090] = 32'hFFFFFFF1;
    // rom_array[28091] = 32'hFFFFFFF1;
    // rom_array[28092] = 32'hFFFFFFF1;
    // rom_array[28093] = 32'hFFFFFFF1;
    // rom_array[28094] = 32'hFFFFFFF1;
    // rom_array[28095] = 32'hFFFFFFF1;
    // rom_array[28096] = 32'hFFFFFFF1;
    // rom_array[28097] = 32'hFFFFFFF1;
    // rom_array[28098] = 32'hFFFFFFF1;
    // rom_array[28099] = 32'hFFFFFFF1;
    // rom_array[28100] = 32'hFFFFFFF1;
    // rom_array[28101] = 32'hFFFFFFF1;
    // rom_array[28102] = 32'hFFFFFFF1;
    // rom_array[28103] = 32'hFFFFFFF1;
    // rom_array[28104] = 32'hFFFFFFF1;
    // rom_array[28105] = 32'hFFFFFFF1;
    // rom_array[28106] = 32'hFFFFFFF1;
    // rom_array[28107] = 32'hFFFFFFF1;
    // rom_array[28108] = 32'hFFFFFFF1;
    // rom_array[28109] = 32'hFFFFFFF0;
    // rom_array[28110] = 32'hFFFFFFF0;
    // rom_array[28111] = 32'hFFFFFFF0;
    // rom_array[28112] = 32'hFFFFFFF0;
    // rom_array[28113] = 32'hFFFFFFF1;
    // rom_array[28114] = 32'hFFFFFFF1;
    // rom_array[28115] = 32'hFFFFFFF1;
    // rom_array[28116] = 32'hFFFFFFF1;
    // rom_array[28117] = 32'hFFFFFFF0;
    // rom_array[28118] = 32'hFFFFFFF0;
    // rom_array[28119] = 32'hFFFFFFF0;
    // rom_array[28120] = 32'hFFFFFFF0;
    // rom_array[28121] = 32'hFFFFFFF1;
    // rom_array[28122] = 32'hFFFFFFF1;
    // rom_array[28123] = 32'hFFFFFFF1;
    // rom_array[28124] = 32'hFFFFFFF1;
    // rom_array[28125] = 32'hFFFFFFF0;
    // rom_array[28126] = 32'hFFFFFFF0;
    // rom_array[28127] = 32'hFFFFFFF0;
    // rom_array[28128] = 32'hFFFFFFF0;
    // rom_array[28129] = 32'hFFFFFFF1;
    // rom_array[28130] = 32'hFFFFFFF1;
    // rom_array[28131] = 32'hFFFFFFF1;
    // rom_array[28132] = 32'hFFFFFFF1;
    // rom_array[28133] = 32'hFFFFFFF0;
    // rom_array[28134] = 32'hFFFFFFF0;
    // rom_array[28135] = 32'hFFFFFFF0;
    // rom_array[28136] = 32'hFFFFFFF0;
    // rom_array[28137] = 32'hFFFFFFF1;
    // rom_array[28138] = 32'hFFFFFFF1;
    // rom_array[28139] = 32'hFFFFFFF1;
    // rom_array[28140] = 32'hFFFFFFF1;
    // rom_array[28141] = 32'hFFFFFFF1;
    // rom_array[28142] = 32'hFFFFFFF1;
    // rom_array[28143] = 32'hFFFFFFF1;
    // rom_array[28144] = 32'hFFFFFFF1;
    // rom_array[28145] = 32'hFFFFFFF1;
    // rom_array[28146] = 32'hFFFFFFF1;
    // rom_array[28147] = 32'hFFFFFFF1;
    // rom_array[28148] = 32'hFFFFFFF1;
    // rom_array[28149] = 32'hFFFFFFF1;
    // rom_array[28150] = 32'hFFFFFFF1;
    // rom_array[28151] = 32'hFFFFFFF1;
    // rom_array[28152] = 32'hFFFFFFF1;
    // rom_array[28153] = 32'hFFFFFFF1;
    // rom_array[28154] = 32'hFFFFFFF1;
    // rom_array[28155] = 32'hFFFFFFF1;
    // rom_array[28156] = 32'hFFFFFFF1;
    // rom_array[28157] = 32'hFFFFFFF1;
    // rom_array[28158] = 32'hFFFFFFF1;
    // rom_array[28159] = 32'hFFFFFFF1;
    // rom_array[28160] = 32'hFFFFFFF1;
    // rom_array[28161] = 32'hFFFFFFF1;
    // rom_array[28162] = 32'hFFFFFFF1;
    // rom_array[28163] = 32'hFFFFFFF1;
    // rom_array[28164] = 32'hFFFFFFF1;
    // rom_array[28165] = 32'hFFFFFFF1;
    // rom_array[28166] = 32'hFFFFFFF1;
    // rom_array[28167] = 32'hFFFFFFF1;
    // rom_array[28168] = 32'hFFFFFFF1;
    // rom_array[28169] = 32'hFFFFFFF1;
    // rom_array[28170] = 32'hFFFFFFF1;
    // rom_array[28171] = 32'hFFFFFFF1;
    // rom_array[28172] = 32'hFFFFFFF1;
    // rom_array[28173] = 32'hFFFFFFF0;
    // rom_array[28174] = 32'hFFFFFFF0;
    // rom_array[28175] = 32'hFFFFFFF0;
    // rom_array[28176] = 32'hFFFFFFF0;
    // rom_array[28177] = 32'hFFFFFFF1;
    // rom_array[28178] = 32'hFFFFFFF1;
    // rom_array[28179] = 32'hFFFFFFF1;
    // rom_array[28180] = 32'hFFFFFFF1;
    // rom_array[28181] = 32'hFFFFFFF0;
    // rom_array[28182] = 32'hFFFFFFF0;
    // rom_array[28183] = 32'hFFFFFFF0;
    // rom_array[28184] = 32'hFFFFFFF0;
    // rom_array[28185] = 32'hFFFFFFF1;
    // rom_array[28186] = 32'hFFFFFFF1;
    // rom_array[28187] = 32'hFFFFFFF1;
    // rom_array[28188] = 32'hFFFFFFF1;
    // rom_array[28189] = 32'hFFFFFFF0;
    // rom_array[28190] = 32'hFFFFFFF0;
    // rom_array[28191] = 32'hFFFFFFF0;
    // rom_array[28192] = 32'hFFFFFFF0;
    // rom_array[28193] = 32'hFFFFFFF1;
    // rom_array[28194] = 32'hFFFFFFF1;
    // rom_array[28195] = 32'hFFFFFFF1;
    // rom_array[28196] = 32'hFFFFFFF1;
    // rom_array[28197] = 32'hFFFFFFF0;
    // rom_array[28198] = 32'hFFFFFFF0;
    // rom_array[28199] = 32'hFFFFFFF0;
    // rom_array[28200] = 32'hFFFFFFF0;
    // rom_array[28201] = 32'hFFFFFFF1;
    // rom_array[28202] = 32'hFFFFFFF1;
    // rom_array[28203] = 32'hFFFFFFF1;
    // rom_array[28204] = 32'hFFFFFFF1;
    // rom_array[28205] = 32'hFFFFFFF0;
    // rom_array[28206] = 32'hFFFFFFF0;
    // rom_array[28207] = 32'hFFFFFFF1;
    // rom_array[28208] = 32'hFFFFFFF1;
    // rom_array[28209] = 32'hFFFFFFF1;
    // rom_array[28210] = 32'hFFFFFFF1;
    // rom_array[28211] = 32'hFFFFFFF1;
    // rom_array[28212] = 32'hFFFFFFF1;
    // rom_array[28213] = 32'hFFFFFFF0;
    // rom_array[28214] = 32'hFFFFFFF0;
    // rom_array[28215] = 32'hFFFFFFF1;
    // rom_array[28216] = 32'hFFFFFFF1;
    // rom_array[28217] = 32'hFFFFFFF1;
    // rom_array[28218] = 32'hFFFFFFF1;
    // rom_array[28219] = 32'hFFFFFFF1;
    // rom_array[28220] = 32'hFFFFFFF1;
    // rom_array[28221] = 32'hFFFFFFF1;
    // rom_array[28222] = 32'hFFFFFFF1;
    // rom_array[28223] = 32'hFFFFFFF1;
    // rom_array[28224] = 32'hFFFFFFF1;
    // rom_array[28225] = 32'hFFFFFFF1;
    // rom_array[28226] = 32'hFFFFFFF1;
    // rom_array[28227] = 32'hFFFFFFF1;
    // rom_array[28228] = 32'hFFFFFFF1;
    // rom_array[28229] = 32'hFFFFFFF1;
    // rom_array[28230] = 32'hFFFFFFF1;
    // rom_array[28231] = 32'hFFFFFFF1;
    // rom_array[28232] = 32'hFFFFFFF1;
    // rom_array[28233] = 32'hFFFFFFF0;
    // rom_array[28234] = 32'hFFFFFFF0;
    // rom_array[28235] = 32'hFFFFFFF1;
    // rom_array[28236] = 32'hFFFFFFF1;
    // rom_array[28237] = 32'hFFFFFFF0;
    // rom_array[28238] = 32'hFFFFFFF0;
    // rom_array[28239] = 32'hFFFFFFF1;
    // rom_array[28240] = 32'hFFFFFFF1;
    // rom_array[28241] = 32'hFFFFFFF0;
    // rom_array[28242] = 32'hFFFFFFF0;
    // rom_array[28243] = 32'hFFFFFFF1;
    // rom_array[28244] = 32'hFFFFFFF1;
    // rom_array[28245] = 32'hFFFFFFF0;
    // rom_array[28246] = 32'hFFFFFFF0;
    // rom_array[28247] = 32'hFFFFFFF1;
    // rom_array[28248] = 32'hFFFFFFF1;
    // rom_array[28249] = 32'hFFFFFFF0;
    // rom_array[28250] = 32'hFFFFFFF0;
    // rom_array[28251] = 32'hFFFFFFF1;
    // rom_array[28252] = 32'hFFFFFFF1;
    // rom_array[28253] = 32'hFFFFFFF0;
    // rom_array[28254] = 32'hFFFFFFF0;
    // rom_array[28255] = 32'hFFFFFFF1;
    // rom_array[28256] = 32'hFFFFFFF1;
    // rom_array[28257] = 32'hFFFFFFF0;
    // rom_array[28258] = 32'hFFFFFFF0;
    // rom_array[28259] = 32'hFFFFFFF1;
    // rom_array[28260] = 32'hFFFFFFF1;
    // rom_array[28261] = 32'hFFFFFFF0;
    // rom_array[28262] = 32'hFFFFFFF0;
    // rom_array[28263] = 32'hFFFFFFF1;
    // rom_array[28264] = 32'hFFFFFFF1;
    // rom_array[28265] = 32'hFFFFFFF0;
    // rom_array[28266] = 32'hFFFFFFF0;
    // rom_array[28267] = 32'hFFFFFFF1;
    // rom_array[28268] = 32'hFFFFFFF1;
    // rom_array[28269] = 32'hFFFFFFF0;
    // rom_array[28270] = 32'hFFFFFFF0;
    // rom_array[28271] = 32'hFFFFFFF1;
    // rom_array[28272] = 32'hFFFFFFF1;
    // rom_array[28273] = 32'hFFFFFFF0;
    // rom_array[28274] = 32'hFFFFFFF0;
    // rom_array[28275] = 32'hFFFFFFF1;
    // rom_array[28276] = 32'hFFFFFFF1;
    // rom_array[28277] = 32'hFFFFFFF0;
    // rom_array[28278] = 32'hFFFFFFF0;
    // rom_array[28279] = 32'hFFFFFFF1;
    // rom_array[28280] = 32'hFFFFFFF1;
    // rom_array[28281] = 32'hFFFFFFF0;
    // rom_array[28282] = 32'hFFFFFFF0;
    // rom_array[28283] = 32'hFFFFFFF0;
    // rom_array[28284] = 32'hFFFFFFF0;
    // rom_array[28285] = 32'hFFFFFFF1;
    // rom_array[28286] = 32'hFFFFFFF1;
    // rom_array[28287] = 32'hFFFFFFF1;
    // rom_array[28288] = 32'hFFFFFFF1;
    // rom_array[28289] = 32'hFFFFFFF0;
    // rom_array[28290] = 32'hFFFFFFF0;
    // rom_array[28291] = 32'hFFFFFFF0;
    // rom_array[28292] = 32'hFFFFFFF0;
    // rom_array[28293] = 32'hFFFFFFF1;
    // rom_array[28294] = 32'hFFFFFFF1;
    // rom_array[28295] = 32'hFFFFFFF1;
    // rom_array[28296] = 32'hFFFFFFF1;
    // rom_array[28297] = 32'hFFFFFFF0;
    // rom_array[28298] = 32'hFFFFFFF0;
    // rom_array[28299] = 32'hFFFFFFF0;
    // rom_array[28300] = 32'hFFFFFFF0;
    // rom_array[28301] = 32'hFFFFFFF1;
    // rom_array[28302] = 32'hFFFFFFF1;
    // rom_array[28303] = 32'hFFFFFFF1;
    // rom_array[28304] = 32'hFFFFFFF1;
    // rom_array[28305] = 32'hFFFFFFF0;
    // rom_array[28306] = 32'hFFFFFFF0;
    // rom_array[28307] = 32'hFFFFFFF0;
    // rom_array[28308] = 32'hFFFFFFF0;
    // rom_array[28309] = 32'hFFFFFFF1;
    // rom_array[28310] = 32'hFFFFFFF1;
    // rom_array[28311] = 32'hFFFFFFF1;
    // rom_array[28312] = 32'hFFFFFFF1;
    // rom_array[28313] = 32'hFFFFFFF0;
    // rom_array[28314] = 32'hFFFFFFF0;
    // rom_array[28315] = 32'hFFFFFFF0;
    // rom_array[28316] = 32'hFFFFFFF0;
    // rom_array[28317] = 32'hFFFFFFF1;
    // rom_array[28318] = 32'hFFFFFFF1;
    // rom_array[28319] = 32'hFFFFFFF1;
    // rom_array[28320] = 32'hFFFFFFF1;
    // rom_array[28321] = 32'hFFFFFFF0;
    // rom_array[28322] = 32'hFFFFFFF0;
    // rom_array[28323] = 32'hFFFFFFF0;
    // rom_array[28324] = 32'hFFFFFFF0;
    // rom_array[28325] = 32'hFFFFFFF1;
    // rom_array[28326] = 32'hFFFFFFF1;
    // rom_array[28327] = 32'hFFFFFFF1;
    // rom_array[28328] = 32'hFFFFFFF1;
    // rom_array[28329] = 32'hFFFFFFF1;
    // rom_array[28330] = 32'hFFFFFFF1;
    // rom_array[28331] = 32'hFFFFFFF1;
    // rom_array[28332] = 32'hFFFFFFF1;
    // rom_array[28333] = 32'hFFFFFFF1;
    // rom_array[28334] = 32'hFFFFFFF1;
    // rom_array[28335] = 32'hFFFFFFF1;
    // rom_array[28336] = 32'hFFFFFFF1;
    // rom_array[28337] = 32'hFFFFFFF1;
    // rom_array[28338] = 32'hFFFFFFF1;
    // rom_array[28339] = 32'hFFFFFFF1;
    // rom_array[28340] = 32'hFFFFFFF1;
    // rom_array[28341] = 32'hFFFFFFF1;
    // rom_array[28342] = 32'hFFFFFFF1;
    // rom_array[28343] = 32'hFFFFFFF1;
    // rom_array[28344] = 32'hFFFFFFF1;
    // rom_array[28345] = 32'hFFFFFFF1;
    // rom_array[28346] = 32'hFFFFFFF1;
    // rom_array[28347] = 32'hFFFFFFF1;
    // rom_array[28348] = 32'hFFFFFFF1;
    // rom_array[28349] = 32'hFFFFFFF1;
    // rom_array[28350] = 32'hFFFFFFF1;
    // rom_array[28351] = 32'hFFFFFFF1;
    // rom_array[28352] = 32'hFFFFFFF1;
    // rom_array[28353] = 32'hFFFFFFF1;
    // rom_array[28354] = 32'hFFFFFFF1;
    // rom_array[28355] = 32'hFFFFFFF1;
    // rom_array[28356] = 32'hFFFFFFF1;
    // rom_array[28357] = 32'hFFFFFFF1;
    // rom_array[28358] = 32'hFFFFFFF1;
    // rom_array[28359] = 32'hFFFFFFF1;
    // rom_array[28360] = 32'hFFFFFFF1;
    // rom_array[28361] = 32'hFFFFFFF1;
    // rom_array[28362] = 32'hFFFFFFF1;
    // rom_array[28363] = 32'hFFFFFFF1;
    // rom_array[28364] = 32'hFFFFFFF1;
    // rom_array[28365] = 32'hFFFFFFF1;
    // rom_array[28366] = 32'hFFFFFFF1;
    // rom_array[28367] = 32'hFFFFFFF1;
    // rom_array[28368] = 32'hFFFFFFF1;
    // rom_array[28369] = 32'hFFFFFFF1;
    // rom_array[28370] = 32'hFFFFFFF1;
    // rom_array[28371] = 32'hFFFFFFF1;
    // rom_array[28372] = 32'hFFFFFFF1;
    // rom_array[28373] = 32'hFFFFFFF1;
    // rom_array[28374] = 32'hFFFFFFF1;
    // rom_array[28375] = 32'hFFFFFFF1;
    // rom_array[28376] = 32'hFFFFFFF1;
    // rom_array[28377] = 32'hFFFFFFF1;
    // rom_array[28378] = 32'hFFFFFFF1;
    // rom_array[28379] = 32'hFFFFFFF1;
    // rom_array[28380] = 32'hFFFFFFF1;
    // rom_array[28381] = 32'hFFFFFFF1;
    // rom_array[28382] = 32'hFFFFFFF1;
    // rom_array[28383] = 32'hFFFFFFF1;
    // rom_array[28384] = 32'hFFFFFFF1;
    // rom_array[28385] = 32'hFFFFFFF1;
    // rom_array[28386] = 32'hFFFFFFF1;
    // rom_array[28387] = 32'hFFFFFFF1;
    // rom_array[28388] = 32'hFFFFFFF1;
    // rom_array[28389] = 32'hFFFFFFF1;
    // rom_array[28390] = 32'hFFFFFFF1;
    // rom_array[28391] = 32'hFFFFFFF1;
    // rom_array[28392] = 32'hFFFFFFF1;
    // rom_array[28393] = 32'hFFFFFFF1;
    // rom_array[28394] = 32'hFFFFFFF1;
    // rom_array[28395] = 32'hFFFFFFF1;
    // rom_array[28396] = 32'hFFFFFFF1;
    // rom_array[28397] = 32'hFFFFFFF1;
    // rom_array[28398] = 32'hFFFFFFF1;
    // rom_array[28399] = 32'hFFFFFFF1;
    // rom_array[28400] = 32'hFFFFFFF1;
    // rom_array[28401] = 32'hFFFFFFF1;
    // rom_array[28402] = 32'hFFFFFFF1;
    // rom_array[28403] = 32'hFFFFFFF1;
    // rom_array[28404] = 32'hFFFFFFF1;
    // rom_array[28405] = 32'hFFFFFFF1;
    // rom_array[28406] = 32'hFFFFFFF1;
    // rom_array[28407] = 32'hFFFFFFF1;
    // rom_array[28408] = 32'hFFFFFFF1;
    // rom_array[28409] = 32'hFFFFFFF1;
    // rom_array[28410] = 32'hFFFFFFF1;
    // rom_array[28411] = 32'hFFFFFFF1;
    // rom_array[28412] = 32'hFFFFFFF1;
    // rom_array[28413] = 32'hFFFFFFF1;
    // rom_array[28414] = 32'hFFFFFFF1;
    // rom_array[28415] = 32'hFFFFFFF1;
    // rom_array[28416] = 32'hFFFFFFF1;
    // rom_array[28417] = 32'hFFFFFFF1;
    // rom_array[28418] = 32'hFFFFFFF1;
    // rom_array[28419] = 32'hFFFFFFF1;
    // rom_array[28420] = 32'hFFFFFFF1;
    // rom_array[28421] = 32'hFFFFFFF1;
    // rom_array[28422] = 32'hFFFFFFF1;
    // rom_array[28423] = 32'hFFFFFFF1;
    // rom_array[28424] = 32'hFFFFFFF1;
    // rom_array[28425] = 32'hFFFFFFF1;
    // rom_array[28426] = 32'hFFFFFFF1;
    // rom_array[28427] = 32'hFFFFFFF1;
    // rom_array[28428] = 32'hFFFFFFF1;
    // rom_array[28429] = 32'hFFFFFFF1;
    // rom_array[28430] = 32'hFFFFFFF1;
    // rom_array[28431] = 32'hFFFFFFF1;
    // rom_array[28432] = 32'hFFFFFFF1;
    // rom_array[28433] = 32'hFFFFFFF1;
    // rom_array[28434] = 32'hFFFFFFF1;
    // rom_array[28435] = 32'hFFFFFFF1;
    // rom_array[28436] = 32'hFFFFFFF1;
    // rom_array[28437] = 32'hFFFFFFF1;
    // rom_array[28438] = 32'hFFFFFFF1;
    // rom_array[28439] = 32'hFFFFFFF1;
    // rom_array[28440] = 32'hFFFFFFF1;
    // rom_array[28441] = 32'hFFFFFFF1;
    // rom_array[28442] = 32'hFFFFFFF1;
    // rom_array[28443] = 32'hFFFFFFF1;
    // rom_array[28444] = 32'hFFFFFFF1;
    // rom_array[28445] = 32'hFFFFFFF1;
    // rom_array[28446] = 32'hFFFFFFF1;
    // rom_array[28447] = 32'hFFFFFFF1;
    // rom_array[28448] = 32'hFFFFFFF1;
    // rom_array[28449] = 32'hFFFFFFF1;
    // rom_array[28450] = 32'hFFFFFFF1;
    // rom_array[28451] = 32'hFFFFFFF1;
    // rom_array[28452] = 32'hFFFFFFF1;
    // rom_array[28453] = 32'hFFFFFFF1;
    // rom_array[28454] = 32'hFFFFFFF1;
    // rom_array[28455] = 32'hFFFFFFF1;
    // rom_array[28456] = 32'hFFFFFFF1;
    // rom_array[28457] = 32'hFFFFFFF1;
    // rom_array[28458] = 32'hFFFFFFF1;
    // rom_array[28459] = 32'hFFFFFFF1;
    // rom_array[28460] = 32'hFFFFFFF1;
    // rom_array[28461] = 32'hFFFFFFF1;
    // rom_array[28462] = 32'hFFFFFFF1;
    // rom_array[28463] = 32'hFFFFFFF1;
    // rom_array[28464] = 32'hFFFFFFF1;
    // rom_array[28465] = 32'hFFFFFFF1;
    // rom_array[28466] = 32'hFFFFFFF1;
    // rom_array[28467] = 32'hFFFFFFF1;
    // rom_array[28468] = 32'hFFFFFFF1;
    // rom_array[28469] = 32'hFFFFFFF1;
    // rom_array[28470] = 32'hFFFFFFF1;
    // rom_array[28471] = 32'hFFFFFFF1;
    // rom_array[28472] = 32'hFFFFFFF1;
    // rom_array[28473] = 32'hFFFFFFF1;
    // rom_array[28474] = 32'hFFFFFFF1;
    // rom_array[28475] = 32'hFFFFFFF1;
    // rom_array[28476] = 32'hFFFFFFF1;
    // rom_array[28477] = 32'hFFFFFFF1;
    // rom_array[28478] = 32'hFFFFFFF1;
    // rom_array[28479] = 32'hFFFFFFF1;
    // rom_array[28480] = 32'hFFFFFFF1;
    // rom_array[28481] = 32'hFFFFFFF1;
    // rom_array[28482] = 32'hFFFFFFF1;
    // rom_array[28483] = 32'hFFFFFFF1;
    // rom_array[28484] = 32'hFFFFFFF1;
    // rom_array[28485] = 32'hFFFFFFF1;
    // rom_array[28486] = 32'hFFFFFFF1;
    // rom_array[28487] = 32'hFFFFFFF1;
    // rom_array[28488] = 32'hFFFFFFF1;
    // rom_array[28489] = 32'hFFFFFFF1;
    // rom_array[28490] = 32'hFFFFFFF1;
    // rom_array[28491] = 32'hFFFFFFF1;
    // rom_array[28492] = 32'hFFFFFFF1;
    // rom_array[28493] = 32'hFFFFFFF1;
    // rom_array[28494] = 32'hFFFFFFF1;
    // rom_array[28495] = 32'hFFFFFFF1;
    // rom_array[28496] = 32'hFFFFFFF1;
    // rom_array[28497] = 32'hFFFFFFF1;
    // rom_array[28498] = 32'hFFFFFFF1;
    // rom_array[28499] = 32'hFFFFFFF1;
    // rom_array[28500] = 32'hFFFFFFF1;
    // rom_array[28501] = 32'hFFFFFFF1;
    // rom_array[28502] = 32'hFFFFFFF1;
    // rom_array[28503] = 32'hFFFFFFF1;
    // rom_array[28504] = 32'hFFFFFFF1;
    // rom_array[28505] = 32'hFFFFFFF1;
    // rom_array[28506] = 32'hFFFFFFF1;
    // rom_array[28507] = 32'hFFFFFFF1;
    // rom_array[28508] = 32'hFFFFFFF1;
    // rom_array[28509] = 32'hFFFFFFF1;
    // rom_array[28510] = 32'hFFFFFFF1;
    // rom_array[28511] = 32'hFFFFFFF1;
    // rom_array[28512] = 32'hFFFFFFF1;
    // rom_array[28513] = 32'hFFFFFFF1;
    // rom_array[28514] = 32'hFFFFFFF1;
    // rom_array[28515] = 32'hFFFFFFF1;
    // rom_array[28516] = 32'hFFFFFFF1;
    // rom_array[28517] = 32'hFFFFFFF1;
    // rom_array[28518] = 32'hFFFFFFF1;
    // rom_array[28519] = 32'hFFFFFFF1;
    // rom_array[28520] = 32'hFFFFFFF1;
    // rom_array[28521] = 32'hFFFFFFF1;
    // rom_array[28522] = 32'hFFFFFFF1;
    // rom_array[28523] = 32'hFFFFFFF1;
    // rom_array[28524] = 32'hFFFFFFF1;
    // rom_array[28525] = 32'hFFFFFFF1;
    // rom_array[28526] = 32'hFFFFFFF1;
    // rom_array[28527] = 32'hFFFFFFF1;
    // rom_array[28528] = 32'hFFFFFFF1;
    // rom_array[28529] = 32'hFFFFFFF1;
    // rom_array[28530] = 32'hFFFFFFF1;
    // rom_array[28531] = 32'hFFFFFFF1;
    // rom_array[28532] = 32'hFFFFFFF1;
    // rom_array[28533] = 32'hFFFFFFF1;
    // rom_array[28534] = 32'hFFFFFFF1;
    // rom_array[28535] = 32'hFFFFFFF1;
    // rom_array[28536] = 32'hFFFFFFF1;
    // rom_array[28537] = 32'hFFFFFFF0;
    // rom_array[28538] = 32'hFFFFFFF0;
    // rom_array[28539] = 32'hFFFFFFF0;
    // rom_array[28540] = 32'hFFFFFFF0;
    // rom_array[28541] = 32'hFFFFFFF1;
    // rom_array[28542] = 32'hFFFFFFF1;
    // rom_array[28543] = 32'hFFFFFFF1;
    // rom_array[28544] = 32'hFFFFFFF1;
    // rom_array[28545] = 32'hFFFFFFF0;
    // rom_array[28546] = 32'hFFFFFFF0;
    // rom_array[28547] = 32'hFFFFFFF0;
    // rom_array[28548] = 32'hFFFFFFF0;
    // rom_array[28549] = 32'hFFFFFFF1;
    // rom_array[28550] = 32'hFFFFFFF1;
    // rom_array[28551] = 32'hFFFFFFF1;
    // rom_array[28552] = 32'hFFFFFFF1;
    // rom_array[28553] = 32'hFFFFFFF0;
    // rom_array[28554] = 32'hFFFFFFF0;
    // rom_array[28555] = 32'hFFFFFFF0;
    // rom_array[28556] = 32'hFFFFFFF0;
    // rom_array[28557] = 32'hFFFFFFF1;
    // rom_array[28558] = 32'hFFFFFFF1;
    // rom_array[28559] = 32'hFFFFFFF1;
    // rom_array[28560] = 32'hFFFFFFF1;
    // rom_array[28561] = 32'hFFFFFFF0;
    // rom_array[28562] = 32'hFFFFFFF0;
    // rom_array[28563] = 32'hFFFFFFF0;
    // rom_array[28564] = 32'hFFFFFFF0;
    // rom_array[28565] = 32'hFFFFFFF1;
    // rom_array[28566] = 32'hFFFFFFF1;
    // rom_array[28567] = 32'hFFFFFFF1;
    // rom_array[28568] = 32'hFFFFFFF1;
    // rom_array[28569] = 32'hFFFFFFF0;
    // rom_array[28570] = 32'hFFFFFFF0;
    // rom_array[28571] = 32'hFFFFFFF0;
    // rom_array[28572] = 32'hFFFFFFF0;
    // rom_array[28573] = 32'hFFFFFFF1;
    // rom_array[28574] = 32'hFFFFFFF1;
    // rom_array[28575] = 32'hFFFFFFF1;
    // rom_array[28576] = 32'hFFFFFFF1;
    // rom_array[28577] = 32'hFFFFFFF0;
    // rom_array[28578] = 32'hFFFFFFF0;
    // rom_array[28579] = 32'hFFFFFFF0;
    // rom_array[28580] = 32'hFFFFFFF0;
    // rom_array[28581] = 32'hFFFFFFF1;
    // rom_array[28582] = 32'hFFFFFFF1;
    // rom_array[28583] = 32'hFFFFFFF1;
    // rom_array[28584] = 32'hFFFFFFF1;
    // rom_array[28585] = 32'hFFFFFFF0;
    // rom_array[28586] = 32'hFFFFFFF0;
    // rom_array[28587] = 32'hFFFFFFF1;
    // rom_array[28588] = 32'hFFFFFFF1;
    // rom_array[28589] = 32'hFFFFFFF0;
    // rom_array[28590] = 32'hFFFFFFF0;
    // rom_array[28591] = 32'hFFFFFFF1;
    // rom_array[28592] = 32'hFFFFFFF1;
    // rom_array[28593] = 32'hFFFFFFF0;
    // rom_array[28594] = 32'hFFFFFFF0;
    // rom_array[28595] = 32'hFFFFFFF1;
    // rom_array[28596] = 32'hFFFFFFF1;
    // rom_array[28597] = 32'hFFFFFFF0;
    // rom_array[28598] = 32'hFFFFFFF0;
    // rom_array[28599] = 32'hFFFFFFF1;
    // rom_array[28600] = 32'hFFFFFFF1;
    // rom_array[28601] = 32'hFFFFFFF0;
    // rom_array[28602] = 32'hFFFFFFF0;
    // rom_array[28603] = 32'hFFFFFFF1;
    // rom_array[28604] = 32'hFFFFFFF1;
    // rom_array[28605] = 32'hFFFFFFF0;
    // rom_array[28606] = 32'hFFFFFFF0;
    // rom_array[28607] = 32'hFFFFFFF1;
    // rom_array[28608] = 32'hFFFFFFF1;
    // rom_array[28609] = 32'hFFFFFFF0;
    // rom_array[28610] = 32'hFFFFFFF0;
    // rom_array[28611] = 32'hFFFFFFF1;
    // rom_array[28612] = 32'hFFFFFFF1;
    // rom_array[28613] = 32'hFFFFFFF0;
    // rom_array[28614] = 32'hFFFFFFF0;
    // rom_array[28615] = 32'hFFFFFFF1;
    // rom_array[28616] = 32'hFFFFFFF1;
    // rom_array[28617] = 32'hFFFFFFF0;
    // rom_array[28618] = 32'hFFFFFFF0;
    // rom_array[28619] = 32'hFFFFFFF0;
    // rom_array[28620] = 32'hFFFFFFF0;
    // rom_array[28621] = 32'hFFFFFFF1;
    // rom_array[28622] = 32'hFFFFFFF1;
    // rom_array[28623] = 32'hFFFFFFF1;
    // rom_array[28624] = 32'hFFFFFFF1;
    // rom_array[28625] = 32'hFFFFFFF0;
    // rom_array[28626] = 32'hFFFFFFF0;
    // rom_array[28627] = 32'hFFFFFFF0;
    // rom_array[28628] = 32'hFFFFFFF0;
    // rom_array[28629] = 32'hFFFFFFF1;
    // rom_array[28630] = 32'hFFFFFFF1;
    // rom_array[28631] = 32'hFFFFFFF1;
    // rom_array[28632] = 32'hFFFFFFF1;
    // rom_array[28633] = 32'hFFFFFFF0;
    // rom_array[28634] = 32'hFFFFFFF0;
    // rom_array[28635] = 32'hFFFFFFF0;
    // rom_array[28636] = 32'hFFFFFFF0;
    // rom_array[28637] = 32'hFFFFFFF1;
    // rom_array[28638] = 32'hFFFFFFF1;
    // rom_array[28639] = 32'hFFFFFFF1;
    // rom_array[28640] = 32'hFFFFFFF1;
    // rom_array[28641] = 32'hFFFFFFF0;
    // rom_array[28642] = 32'hFFFFFFF0;
    // rom_array[28643] = 32'hFFFFFFF0;
    // rom_array[28644] = 32'hFFFFFFF0;
    // rom_array[28645] = 32'hFFFFFFF1;
    // rom_array[28646] = 32'hFFFFFFF1;
    // rom_array[28647] = 32'hFFFFFFF1;
    // rom_array[28648] = 32'hFFFFFFF1;
    // rom_array[28649] = 32'hFFFFFFF0;
    // rom_array[28650] = 32'hFFFFFFF0;
    // rom_array[28651] = 32'hFFFFFFF1;
    // rom_array[28652] = 32'hFFFFFFF1;
    // rom_array[28653] = 32'hFFFFFFF0;
    // rom_array[28654] = 32'hFFFFFFF0;
    // rom_array[28655] = 32'hFFFFFFF1;
    // rom_array[28656] = 32'hFFFFFFF1;
    // rom_array[28657] = 32'hFFFFFFF0;
    // rom_array[28658] = 32'hFFFFFFF0;
    // rom_array[28659] = 32'hFFFFFFF1;
    // rom_array[28660] = 32'hFFFFFFF1;
    // rom_array[28661] = 32'hFFFFFFF0;
    // rom_array[28662] = 32'hFFFFFFF0;
    // rom_array[28663] = 32'hFFFFFFF1;
    // rom_array[28664] = 32'hFFFFFFF1;
    // rom_array[28665] = 32'hFFFFFFF0;
    // rom_array[28666] = 32'hFFFFFFF0;
    // rom_array[28667] = 32'hFFFFFFF1;
    // rom_array[28668] = 32'hFFFFFFF1;
    // rom_array[28669] = 32'hFFFFFFF1;
    // rom_array[28670] = 32'hFFFFFFF1;
    // rom_array[28671] = 32'hFFFFFFF1;
    // rom_array[28672] = 32'hFFFFFFF1;
    // rom_array[28673] = 32'hFFFFFFF0;
    // rom_array[28674] = 32'hFFFFFFF0;
    // rom_array[28675] = 32'hFFFFFFF1;
    // rom_array[28676] = 32'hFFFFFFF1;
    // rom_array[28677] = 32'hFFFFFFF1;
    // rom_array[28678] = 32'hFFFFFFF1;
    // rom_array[28679] = 32'hFFFFFFF1;
    // rom_array[28680] = 32'hFFFFFFF1;
    // rom_array[28681] = 32'hFFFFFFF0;
    // rom_array[28682] = 32'hFFFFFFF0;
    // rom_array[28683] = 32'hFFFFFFF0;
    // rom_array[28684] = 32'hFFFFFFF0;
    // rom_array[28685] = 32'hFFFFFFF1;
    // rom_array[28686] = 32'hFFFFFFF1;
    // rom_array[28687] = 32'hFFFFFFF1;
    // rom_array[28688] = 32'hFFFFFFF1;
    // rom_array[28689] = 32'hFFFFFFF0;
    // rom_array[28690] = 32'hFFFFFFF0;
    // rom_array[28691] = 32'hFFFFFFF0;
    // rom_array[28692] = 32'hFFFFFFF0;
    // rom_array[28693] = 32'hFFFFFFF1;
    // rom_array[28694] = 32'hFFFFFFF1;
    // rom_array[28695] = 32'hFFFFFFF1;
    // rom_array[28696] = 32'hFFFFFFF1;
    // rom_array[28697] = 32'hFFFFFFF1;
    // rom_array[28698] = 32'hFFFFFFF1;
    // rom_array[28699] = 32'hFFFFFFF1;
    // rom_array[28700] = 32'hFFFFFFF1;
    // rom_array[28701] = 32'hFFFFFFF0;
    // rom_array[28702] = 32'hFFFFFFF0;
    // rom_array[28703] = 32'hFFFFFFF0;
    // rom_array[28704] = 32'hFFFFFFF0;
    // rom_array[28705] = 32'hFFFFFFF1;
    // rom_array[28706] = 32'hFFFFFFF1;
    // rom_array[28707] = 32'hFFFFFFF1;
    // rom_array[28708] = 32'hFFFFFFF1;
    // rom_array[28709] = 32'hFFFFFFF0;
    // rom_array[28710] = 32'hFFFFFFF0;
    // rom_array[28711] = 32'hFFFFFFF0;
    // rom_array[28712] = 32'hFFFFFFF0;
    // rom_array[28713] = 32'hFFFFFFF1;
    // rom_array[28714] = 32'hFFFFFFF1;
    // rom_array[28715] = 32'hFFFFFFF1;
    // rom_array[28716] = 32'hFFFFFFF1;
    // rom_array[28717] = 32'hFFFFFFF0;
    // rom_array[28718] = 32'hFFFFFFF0;
    // rom_array[28719] = 32'hFFFFFFF0;
    // rom_array[28720] = 32'hFFFFFFF0;
    // rom_array[28721] = 32'hFFFFFFF1;
    // rom_array[28722] = 32'hFFFFFFF1;
    // rom_array[28723] = 32'hFFFFFFF1;
    // rom_array[28724] = 32'hFFFFFFF1;
    // rom_array[28725] = 32'hFFFFFFF0;
    // rom_array[28726] = 32'hFFFFFFF0;
    // rom_array[28727] = 32'hFFFFFFF0;
    // rom_array[28728] = 32'hFFFFFFF0;
    // rom_array[28729] = 32'hFFFFFFF1;
    // rom_array[28730] = 32'hFFFFFFF1;
    // rom_array[28731] = 32'hFFFFFFF1;
    // rom_array[28732] = 32'hFFFFFFF1;
    // rom_array[28733] = 32'hFFFFFFF0;
    // rom_array[28734] = 32'hFFFFFFF0;
    // rom_array[28735] = 32'hFFFFFFF0;
    // rom_array[28736] = 32'hFFFFFFF0;
    // rom_array[28737] = 32'hFFFFFFF1;
    // rom_array[28738] = 32'hFFFFFFF1;
    // rom_array[28739] = 32'hFFFFFFF1;
    // rom_array[28740] = 32'hFFFFFFF1;
    // rom_array[28741] = 32'hFFFFFFF0;
    // rom_array[28742] = 32'hFFFFFFF0;
    // rom_array[28743] = 32'hFFFFFFF0;
    // rom_array[28744] = 32'hFFFFFFF0;
    // rom_array[28745] = 32'hFFFFFFF1;
    // rom_array[28746] = 32'hFFFFFFF1;
    // rom_array[28747] = 32'hFFFFFFF1;
    // rom_array[28748] = 32'hFFFFFFF1;
    // rom_array[28749] = 32'hFFFFFFF0;
    // rom_array[28750] = 32'hFFFFFFF0;
    // rom_array[28751] = 32'hFFFFFFF0;
    // rom_array[28752] = 32'hFFFFFFF0;
    // rom_array[28753] = 32'hFFFFFFF1;
    // rom_array[28754] = 32'hFFFFFFF1;
    // rom_array[28755] = 32'hFFFFFFF1;
    // rom_array[28756] = 32'hFFFFFFF1;
    // rom_array[28757] = 32'hFFFFFFF0;
    // rom_array[28758] = 32'hFFFFFFF0;
    // rom_array[28759] = 32'hFFFFFFF0;
    // rom_array[28760] = 32'hFFFFFFF0;
    // rom_array[28761] = 32'hFFFFFFF1;
    // rom_array[28762] = 32'hFFFFFFF1;
    // rom_array[28763] = 32'hFFFFFFF1;
    // rom_array[28764] = 32'hFFFFFFF1;
    // rom_array[28765] = 32'hFFFFFFF0;
    // rom_array[28766] = 32'hFFFFFFF0;
    // rom_array[28767] = 32'hFFFFFFF0;
    // rom_array[28768] = 32'hFFFFFFF0;
    // rom_array[28769] = 32'hFFFFFFF1;
    // rom_array[28770] = 32'hFFFFFFF1;
    // rom_array[28771] = 32'hFFFFFFF1;
    // rom_array[28772] = 32'hFFFFFFF1;
    // rom_array[28773] = 32'hFFFFFFF0;
    // rom_array[28774] = 32'hFFFFFFF0;
    // rom_array[28775] = 32'hFFFFFFF0;
    // rom_array[28776] = 32'hFFFFFFF0;
    // rom_array[28777] = 32'hFFFFFFF0;
    // rom_array[28778] = 32'hFFFFFFF0;
    // rom_array[28779] = 32'hFFFFFFF1;
    // rom_array[28780] = 32'hFFFFFFF1;
    // rom_array[28781] = 32'hFFFFFFF0;
    // rom_array[28782] = 32'hFFFFFFF0;
    // rom_array[28783] = 32'hFFFFFFF0;
    // rom_array[28784] = 32'hFFFFFFF0;
    // rom_array[28785] = 32'hFFFFFFF0;
    // rom_array[28786] = 32'hFFFFFFF0;
    // rom_array[28787] = 32'hFFFFFFF1;
    // rom_array[28788] = 32'hFFFFFFF1;
    // rom_array[28789] = 32'hFFFFFFF0;
    // rom_array[28790] = 32'hFFFFFFF0;
    // rom_array[28791] = 32'hFFFFFFF0;
    // rom_array[28792] = 32'hFFFFFFF0;
    // rom_array[28793] = 32'hFFFFFFF1;
    // rom_array[28794] = 32'hFFFFFFF1;
    // rom_array[28795] = 32'hFFFFFFF1;
    // rom_array[28796] = 32'hFFFFFFF1;
    // rom_array[28797] = 32'hFFFFFFF1;
    // rom_array[28798] = 32'hFFFFFFF1;
    // rom_array[28799] = 32'hFFFFFFF1;
    // rom_array[28800] = 32'hFFFFFFF1;
    // rom_array[28801] = 32'hFFFFFFF1;
    // rom_array[28802] = 32'hFFFFFFF1;
    // rom_array[28803] = 32'hFFFFFFF1;
    // rom_array[28804] = 32'hFFFFFFF1;
    // rom_array[28805] = 32'hFFFFFFF1;
    // rom_array[28806] = 32'hFFFFFFF1;
    // rom_array[28807] = 32'hFFFFFFF1;
    // rom_array[28808] = 32'hFFFFFFF1;
    // rom_array[28809] = 32'hFFFFFFF1;
    // rom_array[28810] = 32'hFFFFFFF1;
    // rom_array[28811] = 32'hFFFFFFF1;
    // rom_array[28812] = 32'hFFFFFFF1;
    // rom_array[28813] = 32'hFFFFFFF1;
    // rom_array[28814] = 32'hFFFFFFF1;
    // rom_array[28815] = 32'hFFFFFFF1;
    // rom_array[28816] = 32'hFFFFFFF1;
    // rom_array[28817] = 32'hFFFFFFF1;
    // rom_array[28818] = 32'hFFFFFFF1;
    // rom_array[28819] = 32'hFFFFFFF1;
    // rom_array[28820] = 32'hFFFFFFF1;
    // rom_array[28821] = 32'hFFFFFFF1;
    // rom_array[28822] = 32'hFFFFFFF1;
    // rom_array[28823] = 32'hFFFFFFF1;
    // rom_array[28824] = 32'hFFFFFFF1;
    // rom_array[28825] = 32'hFFFFFFF1;
    // rom_array[28826] = 32'hFFFFFFF1;
    // rom_array[28827] = 32'hFFFFFFF1;
    // rom_array[28828] = 32'hFFFFFFF1;
    // rom_array[28829] = 32'hFFFFFFF0;
    // rom_array[28830] = 32'hFFFFFFF0;
    // rom_array[28831] = 32'hFFFFFFF0;
    // rom_array[28832] = 32'hFFFFFFF0;
    // rom_array[28833] = 32'hFFFFFFF1;
    // rom_array[28834] = 32'hFFFFFFF1;
    // rom_array[28835] = 32'hFFFFFFF1;
    // rom_array[28836] = 32'hFFFFFFF1;
    // rom_array[28837] = 32'hFFFFFFF0;
    // rom_array[28838] = 32'hFFFFFFF0;
    // rom_array[28839] = 32'hFFFFFFF0;
    // rom_array[28840] = 32'hFFFFFFF0;
    // rom_array[28841] = 32'hFFFFFFF1;
    // rom_array[28842] = 32'hFFFFFFF1;
    // rom_array[28843] = 32'hFFFFFFF1;
    // rom_array[28844] = 32'hFFFFFFF1;
    // rom_array[28845] = 32'hFFFFFFF0;
    // rom_array[28846] = 32'hFFFFFFF0;
    // rom_array[28847] = 32'hFFFFFFF0;
    // rom_array[28848] = 32'hFFFFFFF0;
    // rom_array[28849] = 32'hFFFFFFF1;
    // rom_array[28850] = 32'hFFFFFFF1;
    // rom_array[28851] = 32'hFFFFFFF1;
    // rom_array[28852] = 32'hFFFFFFF1;
    // rom_array[28853] = 32'hFFFFFFF0;
    // rom_array[28854] = 32'hFFFFFFF0;
    // rom_array[28855] = 32'hFFFFFFF0;
    // rom_array[28856] = 32'hFFFFFFF0;
    // rom_array[28857] = 32'hFFFFFFF1;
    // rom_array[28858] = 32'hFFFFFFF1;
    // rom_array[28859] = 32'hFFFFFFF1;
    // rom_array[28860] = 32'hFFFFFFF1;
    // rom_array[28861] = 32'hFFFFFFF1;
    // rom_array[28862] = 32'hFFFFFFF1;
    // rom_array[28863] = 32'hFFFFFFF1;
    // rom_array[28864] = 32'hFFFFFFF1;
    // rom_array[28865] = 32'hFFFFFFF1;
    // rom_array[28866] = 32'hFFFFFFF1;
    // rom_array[28867] = 32'hFFFFFFF1;
    // rom_array[28868] = 32'hFFFFFFF1;
    // rom_array[28869] = 32'hFFFFFFF1;
    // rom_array[28870] = 32'hFFFFFFF1;
    // rom_array[28871] = 32'hFFFFFFF1;
    // rom_array[28872] = 32'hFFFFFFF1;
    // rom_array[28873] = 32'hFFFFFFF1;
    // rom_array[28874] = 32'hFFFFFFF1;
    // rom_array[28875] = 32'hFFFFFFF1;
    // rom_array[28876] = 32'hFFFFFFF1;
    // rom_array[28877] = 32'hFFFFFFF0;
    // rom_array[28878] = 32'hFFFFFFF0;
    // rom_array[28879] = 32'hFFFFFFF0;
    // rom_array[28880] = 32'hFFFFFFF0;
    // rom_array[28881] = 32'hFFFFFFF1;
    // rom_array[28882] = 32'hFFFFFFF1;
    // rom_array[28883] = 32'hFFFFFFF1;
    // rom_array[28884] = 32'hFFFFFFF1;
    // rom_array[28885] = 32'hFFFFFFF0;
    // rom_array[28886] = 32'hFFFFFFF0;
    // rom_array[28887] = 32'hFFFFFFF0;
    // rom_array[28888] = 32'hFFFFFFF0;
    // rom_array[28889] = 32'hFFFFFFF1;
    // rom_array[28890] = 32'hFFFFFFF1;
    // rom_array[28891] = 32'hFFFFFFF1;
    // rom_array[28892] = 32'hFFFFFFF1;
    // rom_array[28893] = 32'hFFFFFFF0;
    // rom_array[28894] = 32'hFFFFFFF0;
    // rom_array[28895] = 32'hFFFFFFF0;
    // rom_array[28896] = 32'hFFFFFFF0;
    // rom_array[28897] = 32'hFFFFFFF1;
    // rom_array[28898] = 32'hFFFFFFF1;
    // rom_array[28899] = 32'hFFFFFFF1;
    // rom_array[28900] = 32'hFFFFFFF1;
    // rom_array[28901] = 32'hFFFFFFF0;
    // rom_array[28902] = 32'hFFFFFFF0;
    // rom_array[28903] = 32'hFFFFFFF0;
    // rom_array[28904] = 32'hFFFFFFF0;
    // rom_array[28905] = 32'hFFFFFFF1;
    // rom_array[28906] = 32'hFFFFFFF1;
    // rom_array[28907] = 32'hFFFFFFF1;
    // rom_array[28908] = 32'hFFFFFFF1;
    // rom_array[28909] = 32'hFFFFFFF1;
    // rom_array[28910] = 32'hFFFFFFF1;
    // rom_array[28911] = 32'hFFFFFFF1;
    // rom_array[28912] = 32'hFFFFFFF1;
    // rom_array[28913] = 32'hFFFFFFF1;
    // rom_array[28914] = 32'hFFFFFFF1;
    // rom_array[28915] = 32'hFFFFFFF1;
    // rom_array[28916] = 32'hFFFFFFF1;
    // rom_array[28917] = 32'hFFFFFFF1;
    // rom_array[28918] = 32'hFFFFFFF1;
    // rom_array[28919] = 32'hFFFFFFF1;
    // rom_array[28920] = 32'hFFFFFFF1;
    // rom_array[28921] = 32'hFFFFFFF1;
    // rom_array[28922] = 32'hFFFFFFF1;
    // rom_array[28923] = 32'hFFFFFFF1;
    // rom_array[28924] = 32'hFFFFFFF1;
    // rom_array[28925] = 32'hFFFFFFF1;
    // rom_array[28926] = 32'hFFFFFFF1;
    // rom_array[28927] = 32'hFFFFFFF1;
    // rom_array[28928] = 32'hFFFFFFF1;
    // rom_array[28929] = 32'hFFFFFFF1;
    // rom_array[28930] = 32'hFFFFFFF1;
    // rom_array[28931] = 32'hFFFFFFF1;
    // rom_array[28932] = 32'hFFFFFFF1;
    // rom_array[28933] = 32'hFFFFFFF1;
    // rom_array[28934] = 32'hFFFFFFF1;
    // rom_array[28935] = 32'hFFFFFFF1;
    // rom_array[28936] = 32'hFFFFFFF1;
    // rom_array[28937] = 32'hFFFFFFF1;
    // rom_array[28938] = 32'hFFFFFFF1;
    // rom_array[28939] = 32'hFFFFFFF1;
    // rom_array[28940] = 32'hFFFFFFF1;
    // rom_array[28941] = 32'hFFFFFFF1;
    // rom_array[28942] = 32'hFFFFFFF1;
    // rom_array[28943] = 32'hFFFFFFF1;
    // rom_array[28944] = 32'hFFFFFFF1;
    // rom_array[28945] = 32'hFFFFFFF1;
    // rom_array[28946] = 32'hFFFFFFF1;
    // rom_array[28947] = 32'hFFFFFFF1;
    // rom_array[28948] = 32'hFFFFFFF1;
    // rom_array[28949] = 32'hFFFFFFF1;
    // rom_array[28950] = 32'hFFFFFFF1;
    // rom_array[28951] = 32'hFFFFFFF1;
    // rom_array[28952] = 32'hFFFFFFF1;
    // rom_array[28953] = 32'hFFFFFFF1;
    // rom_array[28954] = 32'hFFFFFFF1;
    // rom_array[28955] = 32'hFFFFFFF1;
    // rom_array[28956] = 32'hFFFFFFF1;
    // rom_array[28957] = 32'hFFFFFFF1;
    // rom_array[28958] = 32'hFFFFFFF1;
    // rom_array[28959] = 32'hFFFFFFF1;
    // rom_array[28960] = 32'hFFFFFFF1;
    // rom_array[28961] = 32'hFFFFFFF1;
    // rom_array[28962] = 32'hFFFFFFF1;
    // rom_array[28963] = 32'hFFFFFFF1;
    // rom_array[28964] = 32'hFFFFFFF1;
    // rom_array[28965] = 32'hFFFFFFF1;
    // rom_array[28966] = 32'hFFFFFFF1;
    // rom_array[28967] = 32'hFFFFFFF1;
    // rom_array[28968] = 32'hFFFFFFF1;
    // rom_array[28969] = 32'hFFFFFFF1;
    // rom_array[28970] = 32'hFFFFFFF1;
    // rom_array[28971] = 32'hFFFFFFF1;
    // rom_array[28972] = 32'hFFFFFFF1;
    // rom_array[28973] = 32'hFFFFFFF0;
    // rom_array[28974] = 32'hFFFFFFF0;
    // rom_array[28975] = 32'hFFFFFFF0;
    // rom_array[28976] = 32'hFFFFFFF0;
    // rom_array[28977] = 32'hFFFFFFF1;
    // rom_array[28978] = 32'hFFFFFFF1;
    // rom_array[28979] = 32'hFFFFFFF1;
    // rom_array[28980] = 32'hFFFFFFF1;
    // rom_array[28981] = 32'hFFFFFFF0;
    // rom_array[28982] = 32'hFFFFFFF0;
    // rom_array[28983] = 32'hFFFFFFF0;
    // rom_array[28984] = 32'hFFFFFFF0;
    // rom_array[28985] = 32'hFFFFFFF1;
    // rom_array[28986] = 32'hFFFFFFF1;
    // rom_array[28987] = 32'hFFFFFFF1;
    // rom_array[28988] = 32'hFFFFFFF1;
    // rom_array[28989] = 32'hFFFFFFF0;
    // rom_array[28990] = 32'hFFFFFFF0;
    // rom_array[28991] = 32'hFFFFFFF0;
    // rom_array[28992] = 32'hFFFFFFF0;
    // rom_array[28993] = 32'hFFFFFFF1;
    // rom_array[28994] = 32'hFFFFFFF1;
    // rom_array[28995] = 32'hFFFFFFF1;
    // rom_array[28996] = 32'hFFFFFFF1;
    // rom_array[28997] = 32'hFFFFFFF0;
    // rom_array[28998] = 32'hFFFFFFF0;
    // rom_array[28999] = 32'hFFFFFFF0;
    // rom_array[29000] = 32'hFFFFFFF0;
    // rom_array[29001] = 32'hFFFFFFF1;
    // rom_array[29002] = 32'hFFFFFFF1;
    // rom_array[29003] = 32'hFFFFFFF1;
    // rom_array[29004] = 32'hFFFFFFF1;
    // rom_array[29005] = 32'hFFFFFFF0;
    // rom_array[29006] = 32'hFFFFFFF0;
    // rom_array[29007] = 32'hFFFFFFF0;
    // rom_array[29008] = 32'hFFFFFFF0;
    // rom_array[29009] = 32'hFFFFFFF1;
    // rom_array[29010] = 32'hFFFFFFF1;
    // rom_array[29011] = 32'hFFFFFFF1;
    // rom_array[29012] = 32'hFFFFFFF1;
    // rom_array[29013] = 32'hFFFFFFF0;
    // rom_array[29014] = 32'hFFFFFFF0;
    // rom_array[29015] = 32'hFFFFFFF0;
    // rom_array[29016] = 32'hFFFFFFF0;
    // rom_array[29017] = 32'hFFFFFFF0;
    // rom_array[29018] = 32'hFFFFFFF0;
    // rom_array[29019] = 32'hFFFFFFF0;
    // rom_array[29020] = 32'hFFFFFFF0;
    // rom_array[29021] = 32'hFFFFFFF1;
    // rom_array[29022] = 32'hFFFFFFF1;
    // rom_array[29023] = 32'hFFFFFFF1;
    // rom_array[29024] = 32'hFFFFFFF1;
    // rom_array[29025] = 32'hFFFFFFF0;
    // rom_array[29026] = 32'hFFFFFFF0;
    // rom_array[29027] = 32'hFFFFFFF0;
    // rom_array[29028] = 32'hFFFFFFF0;
    // rom_array[29029] = 32'hFFFFFFF1;
    // rom_array[29030] = 32'hFFFFFFF1;
    // rom_array[29031] = 32'hFFFFFFF1;
    // rom_array[29032] = 32'hFFFFFFF1;
    // rom_array[29033] = 32'hFFFFFFF0;
    // rom_array[29034] = 32'hFFFFFFF0;
    // rom_array[29035] = 32'hFFFFFFF0;
    // rom_array[29036] = 32'hFFFFFFF0;
    // rom_array[29037] = 32'hFFFFFFF1;
    // rom_array[29038] = 32'hFFFFFFF1;
    // rom_array[29039] = 32'hFFFFFFF1;
    // rom_array[29040] = 32'hFFFFFFF1;
    // rom_array[29041] = 32'hFFFFFFF0;
    // rom_array[29042] = 32'hFFFFFFF0;
    // rom_array[29043] = 32'hFFFFFFF0;
    // rom_array[29044] = 32'hFFFFFFF0;
    // rom_array[29045] = 32'hFFFFFFF1;
    // rom_array[29046] = 32'hFFFFFFF1;
    // rom_array[29047] = 32'hFFFFFFF1;
    // rom_array[29048] = 32'hFFFFFFF1;
    // rom_array[29049] = 32'hFFFFFFF0;
    // rom_array[29050] = 32'hFFFFFFF0;
    // rom_array[29051] = 32'hFFFFFFF0;
    // rom_array[29052] = 32'hFFFFFFF0;
    // rom_array[29053] = 32'hFFFFFFF1;
    // rom_array[29054] = 32'hFFFFFFF1;
    // rom_array[29055] = 32'hFFFFFFF1;
    // rom_array[29056] = 32'hFFFFFFF1;
    // rom_array[29057] = 32'hFFFFFFF0;
    // rom_array[29058] = 32'hFFFFFFF0;
    // rom_array[29059] = 32'hFFFFFFF0;
    // rom_array[29060] = 32'hFFFFFFF0;
    // rom_array[29061] = 32'hFFFFFFF1;
    // rom_array[29062] = 32'hFFFFFFF1;
    // rom_array[29063] = 32'hFFFFFFF1;
    // rom_array[29064] = 32'hFFFFFFF1;
    // rom_array[29065] = 32'hFFFFFFF0;
    // rom_array[29066] = 32'hFFFFFFF0;
    // rom_array[29067] = 32'hFFFFFFF0;
    // rom_array[29068] = 32'hFFFFFFF0;
    // rom_array[29069] = 32'hFFFFFFF1;
    // rom_array[29070] = 32'hFFFFFFF1;
    // rom_array[29071] = 32'hFFFFFFF1;
    // rom_array[29072] = 32'hFFFFFFF1;
    // rom_array[29073] = 32'hFFFFFFF0;
    // rom_array[29074] = 32'hFFFFFFF0;
    // rom_array[29075] = 32'hFFFFFFF0;
    // rom_array[29076] = 32'hFFFFFFF0;
    // rom_array[29077] = 32'hFFFFFFF1;
    // rom_array[29078] = 32'hFFFFFFF1;
    // rom_array[29079] = 32'hFFFFFFF1;
    // rom_array[29080] = 32'hFFFFFFF1;
    // rom_array[29081] = 32'hFFFFFFF0;
    // rom_array[29082] = 32'hFFFFFFF0;
    // rom_array[29083] = 32'hFFFFFFF0;
    // rom_array[29084] = 32'hFFFFFFF0;
    // rom_array[29085] = 32'hFFFFFFF1;
    // rom_array[29086] = 32'hFFFFFFF1;
    // rom_array[29087] = 32'hFFFFFFF1;
    // rom_array[29088] = 32'hFFFFFFF1;
    // rom_array[29089] = 32'hFFFFFFF0;
    // rom_array[29090] = 32'hFFFFFFF0;
    // rom_array[29091] = 32'hFFFFFFF0;
    // rom_array[29092] = 32'hFFFFFFF0;
    // rom_array[29093] = 32'hFFFFFFF1;
    // rom_array[29094] = 32'hFFFFFFF1;
    // rom_array[29095] = 32'hFFFFFFF1;
    // rom_array[29096] = 32'hFFFFFFF1;
    // rom_array[29097] = 32'hFFFFFFF0;
    // rom_array[29098] = 32'hFFFFFFF0;
    // rom_array[29099] = 32'hFFFFFFF0;
    // rom_array[29100] = 32'hFFFFFFF0;
    // rom_array[29101] = 32'hFFFFFFF1;
    // rom_array[29102] = 32'hFFFFFFF1;
    // rom_array[29103] = 32'hFFFFFFF1;
    // rom_array[29104] = 32'hFFFFFFF1;
    // rom_array[29105] = 32'hFFFFFFF0;
    // rom_array[29106] = 32'hFFFFFFF0;
    // rom_array[29107] = 32'hFFFFFFF0;
    // rom_array[29108] = 32'hFFFFFFF0;
    // rom_array[29109] = 32'hFFFFFFF1;
    // rom_array[29110] = 32'hFFFFFFF1;
    // rom_array[29111] = 32'hFFFFFFF1;
    // rom_array[29112] = 32'hFFFFFFF1;
    // rom_array[29113] = 32'hFFFFFFF0;
    // rom_array[29114] = 32'hFFFFFFF0;
    // rom_array[29115] = 32'hFFFFFFF0;
    // rom_array[29116] = 32'hFFFFFFF0;
    // rom_array[29117] = 32'hFFFFFFF1;
    // rom_array[29118] = 32'hFFFFFFF1;
    // rom_array[29119] = 32'hFFFFFFF1;
    // rom_array[29120] = 32'hFFFFFFF1;
    // rom_array[29121] = 32'hFFFFFFF0;
    // rom_array[29122] = 32'hFFFFFFF0;
    // rom_array[29123] = 32'hFFFFFFF0;
    // rom_array[29124] = 32'hFFFFFFF0;
    // rom_array[29125] = 32'hFFFFFFF1;
    // rom_array[29126] = 32'hFFFFFFF1;
    // rom_array[29127] = 32'hFFFFFFF1;
    // rom_array[29128] = 32'hFFFFFFF1;
    // rom_array[29129] = 32'hFFFFFFF0;
    // rom_array[29130] = 32'hFFFFFFF0;
    // rom_array[29131] = 32'hFFFFFFF0;
    // rom_array[29132] = 32'hFFFFFFF0;
    // rom_array[29133] = 32'hFFFFFFF1;
    // rom_array[29134] = 32'hFFFFFFF1;
    // rom_array[29135] = 32'hFFFFFFF1;
    // rom_array[29136] = 32'hFFFFFFF1;
    // rom_array[29137] = 32'hFFFFFFF0;
    // rom_array[29138] = 32'hFFFFFFF0;
    // rom_array[29139] = 32'hFFFFFFF0;
    // rom_array[29140] = 32'hFFFFFFF0;
    // rom_array[29141] = 32'hFFFFFFF1;
    // rom_array[29142] = 32'hFFFFFFF1;
    // rom_array[29143] = 32'hFFFFFFF1;
    // rom_array[29144] = 32'hFFFFFFF1;
    // rom_array[29145] = 32'hFFFFFFF1;
    // rom_array[29146] = 32'hFFFFFFF1;
    // rom_array[29147] = 32'hFFFFFFF1;
    // rom_array[29148] = 32'hFFFFFFF1;
    // rom_array[29149] = 32'hFFFFFFF1;
    // rom_array[29150] = 32'hFFFFFFF1;
    // rom_array[29151] = 32'hFFFFFFF1;
    // rom_array[29152] = 32'hFFFFFFF1;
    // rom_array[29153] = 32'hFFFFFFF1;
    // rom_array[29154] = 32'hFFFFFFF1;
    // rom_array[29155] = 32'hFFFFFFF1;
    // rom_array[29156] = 32'hFFFFFFF1;
    // rom_array[29157] = 32'hFFFFFFF1;
    // rom_array[29158] = 32'hFFFFFFF1;
    // rom_array[29159] = 32'hFFFFFFF1;
    // rom_array[29160] = 32'hFFFFFFF1;
    // rom_array[29161] = 32'hFFFFFFF1;
    // rom_array[29162] = 32'hFFFFFFF1;
    // rom_array[29163] = 32'hFFFFFFF1;
    // rom_array[29164] = 32'hFFFFFFF1;
    // rom_array[29165] = 32'hFFFFFFF1;
    // rom_array[29166] = 32'hFFFFFFF1;
    // rom_array[29167] = 32'hFFFFFFF1;
    // rom_array[29168] = 32'hFFFFFFF1;
    // rom_array[29169] = 32'hFFFFFFF1;
    // rom_array[29170] = 32'hFFFFFFF1;
    // rom_array[29171] = 32'hFFFFFFF1;
    // rom_array[29172] = 32'hFFFFFFF1;
    // rom_array[29173] = 32'hFFFFFFF1;
    // rom_array[29174] = 32'hFFFFFFF1;
    // rom_array[29175] = 32'hFFFFFFF1;
    // rom_array[29176] = 32'hFFFFFFF1;
    // rom_array[29177] = 32'hFFFFFFF1;
    // rom_array[29178] = 32'hFFFFFFF1;
    // rom_array[29179] = 32'hFFFFFFF1;
    // rom_array[29180] = 32'hFFFFFFF1;
    // rom_array[29181] = 32'hFFFFFFF1;
    // rom_array[29182] = 32'hFFFFFFF1;
    // rom_array[29183] = 32'hFFFFFFF1;
    // rom_array[29184] = 32'hFFFFFFF1;
    // rom_array[29185] = 32'hFFFFFFF1;
    // rom_array[29186] = 32'hFFFFFFF1;
    // rom_array[29187] = 32'hFFFFFFF1;
    // rom_array[29188] = 32'hFFFFFFF1;
    // rom_array[29189] = 32'hFFFFFFF1;
    // rom_array[29190] = 32'hFFFFFFF1;
    // rom_array[29191] = 32'hFFFFFFF1;
    // rom_array[29192] = 32'hFFFFFFF1;
    // rom_array[29193] = 32'hFFFFFFF1;
    // rom_array[29194] = 32'hFFFFFFF1;
    // rom_array[29195] = 32'hFFFFFFF1;
    // rom_array[29196] = 32'hFFFFFFF1;
    // rom_array[29197] = 32'hFFFFFFF0;
    // rom_array[29198] = 32'hFFFFFFF0;
    // rom_array[29199] = 32'hFFFFFFF0;
    // rom_array[29200] = 32'hFFFFFFF0;
    // rom_array[29201] = 32'hFFFFFFF1;
    // rom_array[29202] = 32'hFFFFFFF1;
    // rom_array[29203] = 32'hFFFFFFF1;
    // rom_array[29204] = 32'hFFFFFFF1;
    // rom_array[29205] = 32'hFFFFFFF0;
    // rom_array[29206] = 32'hFFFFFFF0;
    // rom_array[29207] = 32'hFFFFFFF0;
    // rom_array[29208] = 32'hFFFFFFF0;
    // rom_array[29209] = 32'hFFFFFFF1;
    // rom_array[29210] = 32'hFFFFFFF1;
    // rom_array[29211] = 32'hFFFFFFF1;
    // rom_array[29212] = 32'hFFFFFFF1;
    // rom_array[29213] = 32'hFFFFFFF0;
    // rom_array[29214] = 32'hFFFFFFF0;
    // rom_array[29215] = 32'hFFFFFFF0;
    // rom_array[29216] = 32'hFFFFFFF0;
    // rom_array[29217] = 32'hFFFFFFF1;
    // rom_array[29218] = 32'hFFFFFFF1;
    // rom_array[29219] = 32'hFFFFFFF1;
    // rom_array[29220] = 32'hFFFFFFF1;
    // rom_array[29221] = 32'hFFFFFFF0;
    // rom_array[29222] = 32'hFFFFFFF0;
    // rom_array[29223] = 32'hFFFFFFF0;
    // rom_array[29224] = 32'hFFFFFFF0;
    // rom_array[29225] = 32'hFFFFFFF1;
    // rom_array[29226] = 32'hFFFFFFF1;
    // rom_array[29227] = 32'hFFFFFFF1;
    // rom_array[29228] = 32'hFFFFFFF1;
    // rom_array[29229] = 32'hFFFFFFF0;
    // rom_array[29230] = 32'hFFFFFFF0;
    // rom_array[29231] = 32'hFFFFFFF0;
    // rom_array[29232] = 32'hFFFFFFF0;
    // rom_array[29233] = 32'hFFFFFFF1;
    // rom_array[29234] = 32'hFFFFFFF1;
    // rom_array[29235] = 32'hFFFFFFF1;
    // rom_array[29236] = 32'hFFFFFFF1;
    // rom_array[29237] = 32'hFFFFFFF0;
    // rom_array[29238] = 32'hFFFFFFF0;
    // rom_array[29239] = 32'hFFFFFFF0;
    // rom_array[29240] = 32'hFFFFFFF0;
    // rom_array[29241] = 32'hFFFFFFF1;
    // rom_array[29242] = 32'hFFFFFFF1;
    // rom_array[29243] = 32'hFFFFFFF1;
    // rom_array[29244] = 32'hFFFFFFF1;
    // rom_array[29245] = 32'hFFFFFFF0;
    // rom_array[29246] = 32'hFFFFFFF0;
    // rom_array[29247] = 32'hFFFFFFF0;
    // rom_array[29248] = 32'hFFFFFFF0;
    // rom_array[29249] = 32'hFFFFFFF1;
    // rom_array[29250] = 32'hFFFFFFF1;
    // rom_array[29251] = 32'hFFFFFFF1;
    // rom_array[29252] = 32'hFFFFFFF1;
    // rom_array[29253] = 32'hFFFFFFF0;
    // rom_array[29254] = 32'hFFFFFFF0;
    // rom_array[29255] = 32'hFFFFFFF0;
    // rom_array[29256] = 32'hFFFFFFF0;
    // rom_array[29257] = 32'hFFFFFFF1;
    // rom_array[29258] = 32'hFFFFFFF1;
    // rom_array[29259] = 32'hFFFFFFF1;
    // rom_array[29260] = 32'hFFFFFFF1;
    // rom_array[29261] = 32'hFFFFFFF0;
    // rom_array[29262] = 32'hFFFFFFF0;
    // rom_array[29263] = 32'hFFFFFFF1;
    // rom_array[29264] = 32'hFFFFFFF1;
    // rom_array[29265] = 32'hFFFFFFF1;
    // rom_array[29266] = 32'hFFFFFFF1;
    // rom_array[29267] = 32'hFFFFFFF1;
    // rom_array[29268] = 32'hFFFFFFF1;
    // rom_array[29269] = 32'hFFFFFFF0;
    // rom_array[29270] = 32'hFFFFFFF0;
    // rom_array[29271] = 32'hFFFFFFF1;
    // rom_array[29272] = 32'hFFFFFFF1;
    // rom_array[29273] = 32'hFFFFFFF1;
    // rom_array[29274] = 32'hFFFFFFF1;
    // rom_array[29275] = 32'hFFFFFFF1;
    // rom_array[29276] = 32'hFFFFFFF1;
    // rom_array[29277] = 32'hFFFFFFF1;
    // rom_array[29278] = 32'hFFFFFFF1;
    // rom_array[29279] = 32'hFFFFFFF1;
    // rom_array[29280] = 32'hFFFFFFF1;
    // rom_array[29281] = 32'hFFFFFFF1;
    // rom_array[29282] = 32'hFFFFFFF1;
    // rom_array[29283] = 32'hFFFFFFF1;
    // rom_array[29284] = 32'hFFFFFFF1;
    // rom_array[29285] = 32'hFFFFFFF1;
    // rom_array[29286] = 32'hFFFFFFF1;
    // rom_array[29287] = 32'hFFFFFFF1;
    // rom_array[29288] = 32'hFFFFFFF1;
    // rom_array[29289] = 32'hFFFFFFF0;
    // rom_array[29290] = 32'hFFFFFFF0;
    // rom_array[29291] = 32'hFFFFFFF1;
    // rom_array[29292] = 32'hFFFFFFF1;
    // rom_array[29293] = 32'hFFFFFFF0;
    // rom_array[29294] = 32'hFFFFFFF0;
    // rom_array[29295] = 32'hFFFFFFF1;
    // rom_array[29296] = 32'hFFFFFFF1;
    // rom_array[29297] = 32'hFFFFFFF0;
    // rom_array[29298] = 32'hFFFFFFF0;
    // rom_array[29299] = 32'hFFFFFFF1;
    // rom_array[29300] = 32'hFFFFFFF1;
    // rom_array[29301] = 32'hFFFFFFF0;
    // rom_array[29302] = 32'hFFFFFFF0;
    // rom_array[29303] = 32'hFFFFFFF1;
    // rom_array[29304] = 32'hFFFFFFF1;
    // rom_array[29305] = 32'hFFFFFFF0;
    // rom_array[29306] = 32'hFFFFFFF0;
    // rom_array[29307] = 32'hFFFFFFF0;
    // rom_array[29308] = 32'hFFFFFFF0;
    // rom_array[29309] = 32'hFFFFFFF1;
    // rom_array[29310] = 32'hFFFFFFF1;
    // rom_array[29311] = 32'hFFFFFFF1;
    // rom_array[29312] = 32'hFFFFFFF1;
    // rom_array[29313] = 32'hFFFFFFF0;
    // rom_array[29314] = 32'hFFFFFFF0;
    // rom_array[29315] = 32'hFFFFFFF0;
    // rom_array[29316] = 32'hFFFFFFF0;
    // rom_array[29317] = 32'hFFFFFFF1;
    // rom_array[29318] = 32'hFFFFFFF1;
    // rom_array[29319] = 32'hFFFFFFF1;
    // rom_array[29320] = 32'hFFFFFFF1;
    // rom_array[29321] = 32'hFFFFFFF0;
    // rom_array[29322] = 32'hFFFFFFF0;
    // rom_array[29323] = 32'hFFFFFFF0;
    // rom_array[29324] = 32'hFFFFFFF0;
    // rom_array[29325] = 32'hFFFFFFF1;
    // rom_array[29326] = 32'hFFFFFFF1;
    // rom_array[29327] = 32'hFFFFFFF1;
    // rom_array[29328] = 32'hFFFFFFF1;
    // rom_array[29329] = 32'hFFFFFFF0;
    // rom_array[29330] = 32'hFFFFFFF0;
    // rom_array[29331] = 32'hFFFFFFF0;
    // rom_array[29332] = 32'hFFFFFFF0;
    // rom_array[29333] = 32'hFFFFFFF1;
    // rom_array[29334] = 32'hFFFFFFF1;
    // rom_array[29335] = 32'hFFFFFFF1;
    // rom_array[29336] = 32'hFFFFFFF1;
    // rom_array[29337] = 32'hFFFFFFF0;
    // rom_array[29338] = 32'hFFFFFFF0;
    // rom_array[29339] = 32'hFFFFFFF0;
    // rom_array[29340] = 32'hFFFFFFF0;
    // rom_array[29341] = 32'hFFFFFFF1;
    // rom_array[29342] = 32'hFFFFFFF1;
    // rom_array[29343] = 32'hFFFFFFF1;
    // rom_array[29344] = 32'hFFFFFFF1;
    // rom_array[29345] = 32'hFFFFFFF0;
    // rom_array[29346] = 32'hFFFFFFF0;
    // rom_array[29347] = 32'hFFFFFFF0;
    // rom_array[29348] = 32'hFFFFFFF0;
    // rom_array[29349] = 32'hFFFFFFF1;
    // rom_array[29350] = 32'hFFFFFFF1;
    // rom_array[29351] = 32'hFFFFFFF1;
    // rom_array[29352] = 32'hFFFFFFF1;
    // rom_array[29353] = 32'hFFFFFFF1;
    // rom_array[29354] = 32'hFFFFFFF1;
    // rom_array[29355] = 32'hFFFFFFF1;
    // rom_array[29356] = 32'hFFFFFFF1;
    // rom_array[29357] = 32'hFFFFFFF1;
    // rom_array[29358] = 32'hFFFFFFF1;
    // rom_array[29359] = 32'hFFFFFFF1;
    // rom_array[29360] = 32'hFFFFFFF1;
    // rom_array[29361] = 32'hFFFFFFF1;
    // rom_array[29362] = 32'hFFFFFFF1;
    // rom_array[29363] = 32'hFFFFFFF1;
    // rom_array[29364] = 32'hFFFFFFF1;
    // rom_array[29365] = 32'hFFFFFFF1;
    // rom_array[29366] = 32'hFFFFFFF1;
    // rom_array[29367] = 32'hFFFFFFF1;
    // rom_array[29368] = 32'hFFFFFFF1;
    // rom_array[29369] = 32'hFFFFFFF1;
    // rom_array[29370] = 32'hFFFFFFF1;
    // rom_array[29371] = 32'hFFFFFFF1;
    // rom_array[29372] = 32'hFFFFFFF1;
    // rom_array[29373] = 32'hFFFFFFF1;
    // rom_array[29374] = 32'hFFFFFFF1;
    // rom_array[29375] = 32'hFFFFFFF1;
    // rom_array[29376] = 32'hFFFFFFF1;
    // rom_array[29377] = 32'hFFFFFFF1;
    // rom_array[29378] = 32'hFFFFFFF1;
    // rom_array[29379] = 32'hFFFFFFF1;
    // rom_array[29380] = 32'hFFFFFFF1;
    // rom_array[29381] = 32'hFFFFFFF1;
    // rom_array[29382] = 32'hFFFFFFF1;
    // rom_array[29383] = 32'hFFFFFFF1;
    // rom_array[29384] = 32'hFFFFFFF1;
    // rom_array[29385] = 32'hFFFFFFF1;
    // rom_array[29386] = 32'hFFFFFFF1;
    // rom_array[29387] = 32'hFFFFFFF1;
    // rom_array[29388] = 32'hFFFFFFF1;
    // rom_array[29389] = 32'hFFFFFFF1;
    // rom_array[29390] = 32'hFFFFFFF1;
    // rom_array[29391] = 32'hFFFFFFF1;
    // rom_array[29392] = 32'hFFFFFFF1;
    // rom_array[29393] = 32'hFFFFFFF1;
    // rom_array[29394] = 32'hFFFFFFF1;
    // rom_array[29395] = 32'hFFFFFFF1;
    // rom_array[29396] = 32'hFFFFFFF1;
    // rom_array[29397] = 32'hFFFFFFF1;
    // rom_array[29398] = 32'hFFFFFFF1;
    // rom_array[29399] = 32'hFFFFFFF1;
    // rom_array[29400] = 32'hFFFFFFF1;
    // rom_array[29401] = 32'hFFFFFFF1;
    // rom_array[29402] = 32'hFFFFFFF1;
    // rom_array[29403] = 32'hFFFFFFF1;
    // rom_array[29404] = 32'hFFFFFFF1;
    // rom_array[29405] = 32'hFFFFFFF1;
    // rom_array[29406] = 32'hFFFFFFF1;
    // rom_array[29407] = 32'hFFFFFFF1;
    // rom_array[29408] = 32'hFFFFFFF1;
    // rom_array[29409] = 32'hFFFFFFF1;
    // rom_array[29410] = 32'hFFFFFFF1;
    // rom_array[29411] = 32'hFFFFFFF1;
    // rom_array[29412] = 32'hFFFFFFF1;
    // rom_array[29413] = 32'hFFFFFFF1;
    // rom_array[29414] = 32'hFFFFFFF1;
    // rom_array[29415] = 32'hFFFFFFF1;
    // rom_array[29416] = 32'hFFFFFFF1;
    // rom_array[29417] = 32'hFFFFFFF1;
    // rom_array[29418] = 32'hFFFFFFF1;
    // rom_array[29419] = 32'hFFFFFFF1;
    // rom_array[29420] = 32'hFFFFFFF1;
    // rom_array[29421] = 32'hFFFFFFF1;
    // rom_array[29422] = 32'hFFFFFFF1;
    // rom_array[29423] = 32'hFFFFFFF1;
    // rom_array[29424] = 32'hFFFFFFF1;
    // rom_array[29425] = 32'hFFFFFFF1;
    // rom_array[29426] = 32'hFFFFFFF1;
    // rom_array[29427] = 32'hFFFFFFF1;
    // rom_array[29428] = 32'hFFFFFFF1;
    // rom_array[29429] = 32'hFFFFFFF1;
    // rom_array[29430] = 32'hFFFFFFF1;
    // rom_array[29431] = 32'hFFFFFFF1;
    // rom_array[29432] = 32'hFFFFFFF1;
    // rom_array[29433] = 32'hFFFFFFF1;
    // rom_array[29434] = 32'hFFFFFFF1;
    // rom_array[29435] = 32'hFFFFFFF1;
    // rom_array[29436] = 32'hFFFFFFF1;
    // rom_array[29437] = 32'hFFFFFFF1;
    // rom_array[29438] = 32'hFFFFFFF1;
    // rom_array[29439] = 32'hFFFFFFF1;
    // rom_array[29440] = 32'hFFFFFFF1;
    // rom_array[29441] = 32'hFFFFFFF1;
    // rom_array[29442] = 32'hFFFFFFF1;
    // rom_array[29443] = 32'hFFFFFFF1;
    // rom_array[29444] = 32'hFFFFFFF1;
    // rom_array[29445] = 32'hFFFFFFF1;
    // rom_array[29446] = 32'hFFFFFFF1;
    // rom_array[29447] = 32'hFFFFFFF1;
    // rom_array[29448] = 32'hFFFFFFF1;
    // rom_array[29449] = 32'hFFFFFFF1;
    // rom_array[29450] = 32'hFFFFFFF1;
    // rom_array[29451] = 32'hFFFFFFF1;
    // rom_array[29452] = 32'hFFFFFFF1;
    // rom_array[29453] = 32'hFFFFFFF1;
    // rom_array[29454] = 32'hFFFFFFF1;
    // rom_array[29455] = 32'hFFFFFFF1;
    // rom_array[29456] = 32'hFFFFFFF1;
    // rom_array[29457] = 32'hFFFFFFF1;
    // rom_array[29458] = 32'hFFFFFFF1;
    // rom_array[29459] = 32'hFFFFFFF1;
    // rom_array[29460] = 32'hFFFFFFF1;
    // rom_array[29461] = 32'hFFFFFFF1;
    // rom_array[29462] = 32'hFFFFFFF1;
    // rom_array[29463] = 32'hFFFFFFF1;
    // rom_array[29464] = 32'hFFFFFFF1;
    // rom_array[29465] = 32'hFFFFFFF1;
    // rom_array[29466] = 32'hFFFFFFF1;
    // rom_array[29467] = 32'hFFFFFFF1;
    // rom_array[29468] = 32'hFFFFFFF1;
    // rom_array[29469] = 32'hFFFFFFF1;
    // rom_array[29470] = 32'hFFFFFFF1;
    // rom_array[29471] = 32'hFFFFFFF1;
    // rom_array[29472] = 32'hFFFFFFF1;
    // rom_array[29473] = 32'hFFFFFFF1;
    // rom_array[29474] = 32'hFFFFFFF1;
    // rom_array[29475] = 32'hFFFFFFF1;
    // rom_array[29476] = 32'hFFFFFFF1;
    // rom_array[29477] = 32'hFFFFFFF1;
    // rom_array[29478] = 32'hFFFFFFF1;
    // rom_array[29479] = 32'hFFFFFFF1;
    // rom_array[29480] = 32'hFFFFFFF1;
    // rom_array[29481] = 32'hFFFFFFF1;
    // rom_array[29482] = 32'hFFFFFFF1;
    // rom_array[29483] = 32'hFFFFFFF1;
    // rom_array[29484] = 32'hFFFFFFF1;
    // rom_array[29485] = 32'hFFFFFFF1;
    // rom_array[29486] = 32'hFFFFFFF1;
    // rom_array[29487] = 32'hFFFFFFF1;
    // rom_array[29488] = 32'hFFFFFFF1;
    // rom_array[29489] = 32'hFFFFFFF1;
    // rom_array[29490] = 32'hFFFFFFF1;
    // rom_array[29491] = 32'hFFFFFFF1;
    // rom_array[29492] = 32'hFFFFFFF1;
    // rom_array[29493] = 32'hFFFFFFF1;
    // rom_array[29494] = 32'hFFFFFFF1;
    // rom_array[29495] = 32'hFFFFFFF1;
    // rom_array[29496] = 32'hFFFFFFF1;
    // rom_array[29497] = 32'hFFFFFFF1;
    // rom_array[29498] = 32'hFFFFFFF1;
    // rom_array[29499] = 32'hFFFFFFF1;
    // rom_array[29500] = 32'hFFFFFFF1;
    // rom_array[29501] = 32'hFFFFFFF1;
    // rom_array[29502] = 32'hFFFFFFF1;
    // rom_array[29503] = 32'hFFFFFFF1;
    // rom_array[29504] = 32'hFFFFFFF1;
    // rom_array[29505] = 32'hFFFFFFF1;
    // rom_array[29506] = 32'hFFFFFFF1;
    // rom_array[29507] = 32'hFFFFFFF1;
    // rom_array[29508] = 32'hFFFFFFF1;
    // rom_array[29509] = 32'hFFFFFFF1;
    // rom_array[29510] = 32'hFFFFFFF1;
    // rom_array[29511] = 32'hFFFFFFF1;
    // rom_array[29512] = 32'hFFFFFFF1;
    // rom_array[29513] = 32'hFFFFFFF1;
    // rom_array[29514] = 32'hFFFFFFF1;
    // rom_array[29515] = 32'hFFFFFFF1;
    // rom_array[29516] = 32'hFFFFFFF1;
    // rom_array[29517] = 32'hFFFFFFF1;
    // rom_array[29518] = 32'hFFFFFFF1;
    // rom_array[29519] = 32'hFFFFFFF1;
    // rom_array[29520] = 32'hFFFFFFF1;
    // rom_array[29521] = 32'hFFFFFFF1;
    // rom_array[29522] = 32'hFFFFFFF1;
    // rom_array[29523] = 32'hFFFFFFF1;
    // rom_array[29524] = 32'hFFFFFFF1;
    // rom_array[29525] = 32'hFFFFFFF1;
    // rom_array[29526] = 32'hFFFFFFF1;
    // rom_array[29527] = 32'hFFFFFFF1;
    // rom_array[29528] = 32'hFFFFFFF1;
    // rom_array[29529] = 32'hFFFFFFF0;
    // rom_array[29530] = 32'hFFFFFFF0;
    // rom_array[29531] = 32'hFFFFFFF1;
    // rom_array[29532] = 32'hFFFFFFF1;
    // rom_array[29533] = 32'hFFFFFFF0;
    // rom_array[29534] = 32'hFFFFFFF0;
    // rom_array[29535] = 32'hFFFFFFF1;
    // rom_array[29536] = 32'hFFFFFFF1;
    // rom_array[29537] = 32'hFFFFFFF0;
    // rom_array[29538] = 32'hFFFFFFF0;
    // rom_array[29539] = 32'hFFFFFFF1;
    // rom_array[29540] = 32'hFFFFFFF1;
    // rom_array[29541] = 32'hFFFFFFF0;
    // rom_array[29542] = 32'hFFFFFFF0;
    // rom_array[29543] = 32'hFFFFFFF1;
    // rom_array[29544] = 32'hFFFFFFF1;
    // rom_array[29545] = 32'hFFFFFFF0;
    // rom_array[29546] = 32'hFFFFFFF0;
    // rom_array[29547] = 32'hFFFFFFF1;
    // rom_array[29548] = 32'hFFFFFFF1;
    // rom_array[29549] = 32'hFFFFFFF0;
    // rom_array[29550] = 32'hFFFFFFF0;
    // rom_array[29551] = 32'hFFFFFFF1;
    // rom_array[29552] = 32'hFFFFFFF1;
    // rom_array[29553] = 32'hFFFFFFF0;
    // rom_array[29554] = 32'hFFFFFFF0;
    // rom_array[29555] = 32'hFFFFFFF1;
    // rom_array[29556] = 32'hFFFFFFF1;
    // rom_array[29557] = 32'hFFFFFFF0;
    // rom_array[29558] = 32'hFFFFFFF0;
    // rom_array[29559] = 32'hFFFFFFF1;
    // rom_array[29560] = 32'hFFFFFFF1;
    // rom_array[29561] = 32'hFFFFFFF0;
    // rom_array[29562] = 32'hFFFFFFF0;
    // rom_array[29563] = 32'hFFFFFFF1;
    // rom_array[29564] = 32'hFFFFFFF1;
    // rom_array[29565] = 32'hFFFFFFF0;
    // rom_array[29566] = 32'hFFFFFFF0;
    // rom_array[29567] = 32'hFFFFFFF1;
    // rom_array[29568] = 32'hFFFFFFF1;
    // rom_array[29569] = 32'hFFFFFFF0;
    // rom_array[29570] = 32'hFFFFFFF0;
    // rom_array[29571] = 32'hFFFFFFF1;
    // rom_array[29572] = 32'hFFFFFFF1;
    // rom_array[29573] = 32'hFFFFFFF0;
    // rom_array[29574] = 32'hFFFFFFF0;
    // rom_array[29575] = 32'hFFFFFFF1;
    // rom_array[29576] = 32'hFFFFFFF1;
    // rom_array[29577] = 32'hFFFFFFF0;
    // rom_array[29578] = 32'hFFFFFFF0;
    // rom_array[29579] = 32'hFFFFFFF1;
    // rom_array[29580] = 32'hFFFFFFF1;
    // rom_array[29581] = 32'hFFFFFFF0;
    // rom_array[29582] = 32'hFFFFFFF0;
    // rom_array[29583] = 32'hFFFFFFF1;
    // rom_array[29584] = 32'hFFFFFFF1;
    // rom_array[29585] = 32'hFFFFFFF0;
    // rom_array[29586] = 32'hFFFFFFF0;
    // rom_array[29587] = 32'hFFFFFFF1;
    // rom_array[29588] = 32'hFFFFFFF1;
    // rom_array[29589] = 32'hFFFFFFF0;
    // rom_array[29590] = 32'hFFFFFFF0;
    // rom_array[29591] = 32'hFFFFFFF1;
    // rom_array[29592] = 32'hFFFFFFF1;
    // rom_array[29593] = 32'hFFFFFFF1;
    // rom_array[29594] = 32'hFFFFFFF1;
    // rom_array[29595] = 32'hFFFFFFF1;
    // rom_array[29596] = 32'hFFFFFFF1;
    // rom_array[29597] = 32'hFFFFFFF1;
    // rom_array[29598] = 32'hFFFFFFF1;
    // rom_array[29599] = 32'hFFFFFFF1;
    // rom_array[29600] = 32'hFFFFFFF1;
    // rom_array[29601] = 32'hFFFFFFF1;
    // rom_array[29602] = 32'hFFFFFFF1;
    // rom_array[29603] = 32'hFFFFFFF1;
    // rom_array[29604] = 32'hFFFFFFF1;
    // rom_array[29605] = 32'hFFFFFFF1;
    // rom_array[29606] = 32'hFFFFFFF1;
    // rom_array[29607] = 32'hFFFFFFF1;
    // rom_array[29608] = 32'hFFFFFFF1;
    // rom_array[29609] = 32'hFFFFFFF1;
    // rom_array[29610] = 32'hFFFFFFF1;
    // rom_array[29611] = 32'hFFFFFFF1;
    // rom_array[29612] = 32'hFFFFFFF1;
    // rom_array[29613] = 32'hFFFFFFF1;
    // rom_array[29614] = 32'hFFFFFFF1;
    // rom_array[29615] = 32'hFFFFFFF1;
    // rom_array[29616] = 32'hFFFFFFF1;
    // rom_array[29617] = 32'hFFFFFFF1;
    // rom_array[29618] = 32'hFFFFFFF1;
    // rom_array[29619] = 32'hFFFFFFF1;
    // rom_array[29620] = 32'hFFFFFFF1;
    // rom_array[29621] = 32'hFFFFFFF1;
    // rom_array[29622] = 32'hFFFFFFF1;
    // rom_array[29623] = 32'hFFFFFFF1;
    // rom_array[29624] = 32'hFFFFFFF1;
    // rom_array[29625] = 32'hFFFFFFF1;
    // rom_array[29626] = 32'hFFFFFFF1;
    // rom_array[29627] = 32'hFFFFFFF1;
    // rom_array[29628] = 32'hFFFFFFF1;
    // rom_array[29629] = 32'hFFFFFFF1;
    // rom_array[29630] = 32'hFFFFFFF1;
    // rom_array[29631] = 32'hFFFFFFF1;
    // rom_array[29632] = 32'hFFFFFFF1;
    // rom_array[29633] = 32'hFFFFFFF1;
    // rom_array[29634] = 32'hFFFFFFF1;
    // rom_array[29635] = 32'hFFFFFFF1;
    // rom_array[29636] = 32'hFFFFFFF1;
    // rom_array[29637] = 32'hFFFFFFF1;
    // rom_array[29638] = 32'hFFFFFFF1;
    // rom_array[29639] = 32'hFFFFFFF1;
    // rom_array[29640] = 32'hFFFFFFF1;
    // rom_array[29641] = 32'hFFFFFFF1;
    // rom_array[29642] = 32'hFFFFFFF1;
    // rom_array[29643] = 32'hFFFFFFF1;
    // rom_array[29644] = 32'hFFFFFFF1;
    // rom_array[29645] = 32'hFFFFFFF1;
    // rom_array[29646] = 32'hFFFFFFF1;
    // rom_array[29647] = 32'hFFFFFFF1;
    // rom_array[29648] = 32'hFFFFFFF1;
    // rom_array[29649] = 32'hFFFFFFF1;
    // rom_array[29650] = 32'hFFFFFFF1;
    // rom_array[29651] = 32'hFFFFFFF1;
    // rom_array[29652] = 32'hFFFFFFF1;
    // rom_array[29653] = 32'hFFFFFFF1;
    // rom_array[29654] = 32'hFFFFFFF1;
    // rom_array[29655] = 32'hFFFFFFF1;
    // rom_array[29656] = 32'hFFFFFFF1;
    // rom_array[29657] = 32'hFFFFFFF0;
    // rom_array[29658] = 32'hFFFFFFF0;
    // rom_array[29659] = 32'hFFFFFFF1;
    // rom_array[29660] = 32'hFFFFFFF1;
    // rom_array[29661] = 32'hFFFFFFF0;
    // rom_array[29662] = 32'hFFFFFFF0;
    // rom_array[29663] = 32'hFFFFFFF1;
    // rom_array[29664] = 32'hFFFFFFF1;
    // rom_array[29665] = 32'hFFFFFFF0;
    // rom_array[29666] = 32'hFFFFFFF0;
    // rom_array[29667] = 32'hFFFFFFF1;
    // rom_array[29668] = 32'hFFFFFFF1;
    // rom_array[29669] = 32'hFFFFFFF0;
    // rom_array[29670] = 32'hFFFFFFF0;
    // rom_array[29671] = 32'hFFFFFFF1;
    // rom_array[29672] = 32'hFFFFFFF1;
    // rom_array[29673] = 32'hFFFFFFF0;
    // rom_array[29674] = 32'hFFFFFFF0;
    // rom_array[29675] = 32'hFFFFFFF1;
    // rom_array[29676] = 32'hFFFFFFF1;
    // rom_array[29677] = 32'hFFFFFFF0;
    // rom_array[29678] = 32'hFFFFFFF0;
    // rom_array[29679] = 32'hFFFFFFF1;
    // rom_array[29680] = 32'hFFFFFFF1;
    // rom_array[29681] = 32'hFFFFFFF0;
    // rom_array[29682] = 32'hFFFFFFF0;
    // rom_array[29683] = 32'hFFFFFFF1;
    // rom_array[29684] = 32'hFFFFFFF1;
    // rom_array[29685] = 32'hFFFFFFF0;
    // rom_array[29686] = 32'hFFFFFFF0;
    // rom_array[29687] = 32'hFFFFFFF1;
    // rom_array[29688] = 32'hFFFFFFF1;
    // rom_array[29689] = 32'hFFFFFFF0;
    // rom_array[29690] = 32'hFFFFFFF0;
    // rom_array[29691] = 32'hFFFFFFF1;
    // rom_array[29692] = 32'hFFFFFFF1;
    // rom_array[29693] = 32'hFFFFFFF0;
    // rom_array[29694] = 32'hFFFFFFF0;
    // rom_array[29695] = 32'hFFFFFFF1;
    // rom_array[29696] = 32'hFFFFFFF1;
    // rom_array[29697] = 32'hFFFFFFF0;
    // rom_array[29698] = 32'hFFFFFFF0;
    // rom_array[29699] = 32'hFFFFFFF1;
    // rom_array[29700] = 32'hFFFFFFF1;
    // rom_array[29701] = 32'hFFFFFFF0;
    // rom_array[29702] = 32'hFFFFFFF0;
    // rom_array[29703] = 32'hFFFFFFF1;
    // rom_array[29704] = 32'hFFFFFFF1;
    // rom_array[29705] = 32'hFFFFFFF0;
    // rom_array[29706] = 32'hFFFFFFF0;
    // rom_array[29707] = 32'hFFFFFFF1;
    // rom_array[29708] = 32'hFFFFFFF1;
    // rom_array[29709] = 32'hFFFFFFF0;
    // rom_array[29710] = 32'hFFFFFFF0;
    // rom_array[29711] = 32'hFFFFFFF1;
    // rom_array[29712] = 32'hFFFFFFF1;
    // rom_array[29713] = 32'hFFFFFFF0;
    // rom_array[29714] = 32'hFFFFFFF0;
    // rom_array[29715] = 32'hFFFFFFF1;
    // rom_array[29716] = 32'hFFFFFFF1;
    // rom_array[29717] = 32'hFFFFFFF0;
    // rom_array[29718] = 32'hFFFFFFF0;
    // rom_array[29719] = 32'hFFFFFFF1;
    // rom_array[29720] = 32'hFFFFFFF1;
    // rom_array[29721] = 32'hFFFFFFF1;
    // rom_array[29722] = 32'hFFFFFFF1;
    // rom_array[29723] = 32'hFFFFFFF1;
    // rom_array[29724] = 32'hFFFFFFF1;
    // rom_array[29725] = 32'hFFFFFFF1;
    // rom_array[29726] = 32'hFFFFFFF1;
    // rom_array[29727] = 32'hFFFFFFF1;
    // rom_array[29728] = 32'hFFFFFFF1;
    // rom_array[29729] = 32'hFFFFFFF1;
    // rom_array[29730] = 32'hFFFFFFF1;
    // rom_array[29731] = 32'hFFFFFFF1;
    // rom_array[29732] = 32'hFFFFFFF1;
    // rom_array[29733] = 32'hFFFFFFF1;
    // rom_array[29734] = 32'hFFFFFFF1;
    // rom_array[29735] = 32'hFFFFFFF1;
    // rom_array[29736] = 32'hFFFFFFF1;
    // rom_array[29737] = 32'hFFFFFFF1;
    // rom_array[29738] = 32'hFFFFFFF1;
    // rom_array[29739] = 32'hFFFFFFF1;
    // rom_array[29740] = 32'hFFFFFFF1;
    // rom_array[29741] = 32'hFFFFFFF1;
    // rom_array[29742] = 32'hFFFFFFF1;
    // rom_array[29743] = 32'hFFFFFFF1;
    // rom_array[29744] = 32'hFFFFFFF1;
    // rom_array[29745] = 32'hFFFFFFF1;
    // rom_array[29746] = 32'hFFFFFFF1;
    // rom_array[29747] = 32'hFFFFFFF1;
    // rom_array[29748] = 32'hFFFFFFF1;
    // rom_array[29749] = 32'hFFFFFFF1;
    // rom_array[29750] = 32'hFFFFFFF1;
    // rom_array[29751] = 32'hFFFFFFF1;
    // rom_array[29752] = 32'hFFFFFFF1;
    // rom_array[29753] = 32'hFFFFFFF1;
    // rom_array[29754] = 32'hFFFFFFF1;
    // rom_array[29755] = 32'hFFFFFFF1;
    // rom_array[29756] = 32'hFFFFFFF1;
    // rom_array[29757] = 32'hFFFFFFF1;
    // rom_array[29758] = 32'hFFFFFFF1;
    // rom_array[29759] = 32'hFFFFFFF1;
    // rom_array[29760] = 32'hFFFFFFF1;
    // rom_array[29761] = 32'hFFFFFFF1;
    // rom_array[29762] = 32'hFFFFFFF1;
    // rom_array[29763] = 32'hFFFFFFF1;
    // rom_array[29764] = 32'hFFFFFFF1;
    // rom_array[29765] = 32'hFFFFFFF1;
    // rom_array[29766] = 32'hFFFFFFF1;
    // rom_array[29767] = 32'hFFFFFFF1;
    // rom_array[29768] = 32'hFFFFFFF1;
    // rom_array[29769] = 32'hFFFFFFF1;
    // rom_array[29770] = 32'hFFFFFFF1;
    // rom_array[29771] = 32'hFFFFFFF1;
    // rom_array[29772] = 32'hFFFFFFF1;
    // rom_array[29773] = 32'hFFFFFFF1;
    // rom_array[29774] = 32'hFFFFFFF1;
    // rom_array[29775] = 32'hFFFFFFF1;
    // rom_array[29776] = 32'hFFFFFFF1;
    // rom_array[29777] = 32'hFFFFFFF1;
    // rom_array[29778] = 32'hFFFFFFF1;
    // rom_array[29779] = 32'hFFFFFFF1;
    // rom_array[29780] = 32'hFFFFFFF1;
    // rom_array[29781] = 32'hFFFFFFF1;
    // rom_array[29782] = 32'hFFFFFFF1;
    // rom_array[29783] = 32'hFFFFFFF1;
    // rom_array[29784] = 32'hFFFFFFF1;
    // rom_array[29785] = 32'hFFFFFFF1;
    // rom_array[29786] = 32'hFFFFFFF1;
    // rom_array[29787] = 32'hFFFFFFF1;
    // rom_array[29788] = 32'hFFFFFFF1;
    // rom_array[29789] = 32'hFFFFFFF1;
    // rom_array[29790] = 32'hFFFFFFF1;
    // rom_array[29791] = 32'hFFFFFFF1;
    // rom_array[29792] = 32'hFFFFFFF1;
    // rom_array[29793] = 32'hFFFFFFF1;
    // rom_array[29794] = 32'hFFFFFFF1;
    // rom_array[29795] = 32'hFFFFFFF1;
    // rom_array[29796] = 32'hFFFFFFF1;
    // rom_array[29797] = 32'hFFFFFFF1;
    // rom_array[29798] = 32'hFFFFFFF1;
    // rom_array[29799] = 32'hFFFFFFF1;
    // rom_array[29800] = 32'hFFFFFFF1;
    // rom_array[29801] = 32'hFFFFFFF1;
    // rom_array[29802] = 32'hFFFFFFF1;
    // rom_array[29803] = 32'hFFFFFFF1;
    // rom_array[29804] = 32'hFFFFFFF1;
    // rom_array[29805] = 32'hFFFFFFF1;
    // rom_array[29806] = 32'hFFFFFFF1;
    // rom_array[29807] = 32'hFFFFFFF1;
    // rom_array[29808] = 32'hFFFFFFF1;
    // rom_array[29809] = 32'hFFFFFFF1;
    // rom_array[29810] = 32'hFFFFFFF1;
    // rom_array[29811] = 32'hFFFFFFF1;
    // rom_array[29812] = 32'hFFFFFFF1;
    // rom_array[29813] = 32'hFFFFFFF1;
    // rom_array[29814] = 32'hFFFFFFF1;
    // rom_array[29815] = 32'hFFFFFFF1;
    // rom_array[29816] = 32'hFFFFFFF1;
    // rom_array[29817] = 32'hFFFFFFF1;
    // rom_array[29818] = 32'hFFFFFFF1;
    // rom_array[29819] = 32'hFFFFFFF1;
    // rom_array[29820] = 32'hFFFFFFF1;
    // rom_array[29821] = 32'hFFFFFFF1;
    // rom_array[29822] = 32'hFFFFFFF1;
    // rom_array[29823] = 32'hFFFFFFF1;
    // rom_array[29824] = 32'hFFFFFFF1;
    // rom_array[29825] = 32'hFFFFFFF1;
    // rom_array[29826] = 32'hFFFFFFF1;
    // rom_array[29827] = 32'hFFFFFFF1;
    // rom_array[29828] = 32'hFFFFFFF1;
    // rom_array[29829] = 32'hFFFFFFF1;
    // rom_array[29830] = 32'hFFFFFFF1;
    // rom_array[29831] = 32'hFFFFFFF1;
    // rom_array[29832] = 32'hFFFFFFF1;
    // rom_array[29833] = 32'hFFFFFFF1;
    // rom_array[29834] = 32'hFFFFFFF1;
    // rom_array[29835] = 32'hFFFFFFF1;
    // rom_array[29836] = 32'hFFFFFFF1;
    // rom_array[29837] = 32'hFFFFFFF1;
    // rom_array[29838] = 32'hFFFFFFF1;
    // rom_array[29839] = 32'hFFFFFFF1;
    // rom_array[29840] = 32'hFFFFFFF1;
    // rom_array[29841] = 32'hFFFFFFF1;
    // rom_array[29842] = 32'hFFFFFFF1;
    // rom_array[29843] = 32'hFFFFFFF1;
    // rom_array[29844] = 32'hFFFFFFF1;
    // rom_array[29845] = 32'hFFFFFFF1;
    // rom_array[29846] = 32'hFFFFFFF1;
    // rom_array[29847] = 32'hFFFFFFF1;
    // rom_array[29848] = 32'hFFFFFFF1;
    // rom_array[29849] = 32'hFFFFFFF0;
    // rom_array[29850] = 32'hFFFFFFF0;
    // rom_array[29851] = 32'hFFFFFFF1;
    // rom_array[29852] = 32'hFFFFFFF1;
    // rom_array[29853] = 32'hFFFFFFF0;
    // rom_array[29854] = 32'hFFFFFFF0;
    // rom_array[29855] = 32'hFFFFFFF0;
    // rom_array[29856] = 32'hFFFFFFF0;
    // rom_array[29857] = 32'hFFFFFFF0;
    // rom_array[29858] = 32'hFFFFFFF0;
    // rom_array[29859] = 32'hFFFFFFF1;
    // rom_array[29860] = 32'hFFFFFFF1;
    // rom_array[29861] = 32'hFFFFFFF0;
    // rom_array[29862] = 32'hFFFFFFF0;
    // rom_array[29863] = 32'hFFFFFFF0;
    // rom_array[29864] = 32'hFFFFFFF0;
    // rom_array[29865] = 32'hFFFFFFF1;
    // rom_array[29866] = 32'hFFFFFFF1;
    // rom_array[29867] = 32'hFFFFFFF1;
    // rom_array[29868] = 32'hFFFFFFF1;
    // rom_array[29869] = 32'hFFFFFFF0;
    // rom_array[29870] = 32'hFFFFFFF0;
    // rom_array[29871] = 32'hFFFFFFF0;
    // rom_array[29872] = 32'hFFFFFFF0;
    // rom_array[29873] = 32'hFFFFFFF1;
    // rom_array[29874] = 32'hFFFFFFF1;
    // rom_array[29875] = 32'hFFFFFFF1;
    // rom_array[29876] = 32'hFFFFFFF1;
    // rom_array[29877] = 32'hFFFFFFF0;
    // rom_array[29878] = 32'hFFFFFFF0;
    // rom_array[29879] = 32'hFFFFFFF0;
    // rom_array[29880] = 32'hFFFFFFF0;
    // rom_array[29881] = 32'hFFFFFFF1;
    // rom_array[29882] = 32'hFFFFFFF1;
    // rom_array[29883] = 32'hFFFFFFF1;
    // rom_array[29884] = 32'hFFFFFFF1;
    // rom_array[29885] = 32'hFFFFFFF0;
    // rom_array[29886] = 32'hFFFFFFF0;
    // rom_array[29887] = 32'hFFFFFFF0;
    // rom_array[29888] = 32'hFFFFFFF0;
    // rom_array[29889] = 32'hFFFFFFF1;
    // rom_array[29890] = 32'hFFFFFFF1;
    // rom_array[29891] = 32'hFFFFFFF1;
    // rom_array[29892] = 32'hFFFFFFF1;
    // rom_array[29893] = 32'hFFFFFFF0;
    // rom_array[29894] = 32'hFFFFFFF0;
    // rom_array[29895] = 32'hFFFFFFF0;
    // rom_array[29896] = 32'hFFFFFFF0;
    // rom_array[29897] = 32'hFFFFFFF1;
    // rom_array[29898] = 32'hFFFFFFF1;
    // rom_array[29899] = 32'hFFFFFFF1;
    // rom_array[29900] = 32'hFFFFFFF1;
    // rom_array[29901] = 32'hFFFFFFF0;
    // rom_array[29902] = 32'hFFFFFFF0;
    // rom_array[29903] = 32'hFFFFFFF0;
    // rom_array[29904] = 32'hFFFFFFF0;
    // rom_array[29905] = 32'hFFFFFFF1;
    // rom_array[29906] = 32'hFFFFFFF1;
    // rom_array[29907] = 32'hFFFFFFF1;
    // rom_array[29908] = 32'hFFFFFFF1;
    // rom_array[29909] = 32'hFFFFFFF0;
    // rom_array[29910] = 32'hFFFFFFF0;
    // rom_array[29911] = 32'hFFFFFFF0;
    // rom_array[29912] = 32'hFFFFFFF0;
    // rom_array[29913] = 32'hFFFFFFF1;
    // rom_array[29914] = 32'hFFFFFFF1;
    // rom_array[29915] = 32'hFFFFFFF1;
    // rom_array[29916] = 32'hFFFFFFF1;
    // rom_array[29917] = 32'hFFFFFFF0;
    // rom_array[29918] = 32'hFFFFFFF0;
    // rom_array[29919] = 32'hFFFFFFF0;
    // rom_array[29920] = 32'hFFFFFFF0;
    // rom_array[29921] = 32'hFFFFFFF1;
    // rom_array[29922] = 32'hFFFFFFF1;
    // rom_array[29923] = 32'hFFFFFFF1;
    // rom_array[29924] = 32'hFFFFFFF1;
    // rom_array[29925] = 32'hFFFFFFF0;
    // rom_array[29926] = 32'hFFFFFFF0;
    // rom_array[29927] = 32'hFFFFFFF0;
    // rom_array[29928] = 32'hFFFFFFF0;
    // rom_array[29929] = 32'hFFFFFFF0;
    // rom_array[29930] = 32'hFFFFFFF0;
    // rom_array[29931] = 32'hFFFFFFF1;
    // rom_array[29932] = 32'hFFFFFFF1;
    // rom_array[29933] = 32'hFFFFFFF0;
    // rom_array[29934] = 32'hFFFFFFF0;
    // rom_array[29935] = 32'hFFFFFFF0;
    // rom_array[29936] = 32'hFFFFFFF0;
    // rom_array[29937] = 32'hFFFFFFF0;
    // rom_array[29938] = 32'hFFFFFFF0;
    // rom_array[29939] = 32'hFFFFFFF1;
    // rom_array[29940] = 32'hFFFFFFF1;
    // rom_array[29941] = 32'hFFFFFFF0;
    // rom_array[29942] = 32'hFFFFFFF0;
    // rom_array[29943] = 32'hFFFFFFF0;
    // rom_array[29944] = 32'hFFFFFFF0;
    // rom_array[29945] = 32'hFFFFFFF1;
    // rom_array[29946] = 32'hFFFFFFF1;
    // rom_array[29947] = 32'hFFFFFFF1;
    // rom_array[29948] = 32'hFFFFFFF1;
    // rom_array[29949] = 32'hFFFFFFF0;
    // rom_array[29950] = 32'hFFFFFFF0;
    // rom_array[29951] = 32'hFFFFFFF0;
    // rom_array[29952] = 32'hFFFFFFF0;
    // rom_array[29953] = 32'hFFFFFFF1;
    // rom_array[29954] = 32'hFFFFFFF1;
    // rom_array[29955] = 32'hFFFFFFF1;
    // rom_array[29956] = 32'hFFFFFFF1;
    // rom_array[29957] = 32'hFFFFFFF0;
    // rom_array[29958] = 32'hFFFFFFF0;
    // rom_array[29959] = 32'hFFFFFFF0;
    // rom_array[29960] = 32'hFFFFFFF0;
    // rom_array[29961] = 32'hFFFFFFF1;
    // rom_array[29962] = 32'hFFFFFFF1;
    // rom_array[29963] = 32'hFFFFFFF1;
    // rom_array[29964] = 32'hFFFFFFF1;
    // rom_array[29965] = 32'hFFFFFFF0;
    // rom_array[29966] = 32'hFFFFFFF0;
    // rom_array[29967] = 32'hFFFFFFF0;
    // rom_array[29968] = 32'hFFFFFFF0;
    // rom_array[29969] = 32'hFFFFFFF1;
    // rom_array[29970] = 32'hFFFFFFF1;
    // rom_array[29971] = 32'hFFFFFFF1;
    // rom_array[29972] = 32'hFFFFFFF1;
    // rom_array[29973] = 32'hFFFFFFF0;
    // rom_array[29974] = 32'hFFFFFFF0;
    // rom_array[29975] = 32'hFFFFFFF0;
    // rom_array[29976] = 32'hFFFFFFF0;
    // rom_array[29977] = 32'hFFFFFFF0;
    // rom_array[29978] = 32'hFFFFFFF0;
    // rom_array[29979] = 32'hFFFFFFF0;
    // rom_array[29980] = 32'hFFFFFFF0;
    // rom_array[29981] = 32'hFFFFFFF0;
    // rom_array[29982] = 32'hFFFFFFF0;
    // rom_array[29983] = 32'hFFFFFFF1;
    // rom_array[29984] = 32'hFFFFFFF1;
    // rom_array[29985] = 32'hFFFFFFF0;
    // rom_array[29986] = 32'hFFFFFFF0;
    // rom_array[29987] = 32'hFFFFFFF0;
    // rom_array[29988] = 32'hFFFFFFF0;
    // rom_array[29989] = 32'hFFFFFFF0;
    // rom_array[29990] = 32'hFFFFFFF0;
    // rom_array[29991] = 32'hFFFFFFF1;
    // rom_array[29992] = 32'hFFFFFFF1;
    // rom_array[29993] = 32'hFFFFFFF0;
    // rom_array[29994] = 32'hFFFFFFF0;
    // rom_array[29995] = 32'hFFFFFFF0;
    // rom_array[29996] = 32'hFFFFFFF0;
    // rom_array[29997] = 32'hFFFFFFF1;
    // rom_array[29998] = 32'hFFFFFFF1;
    // rom_array[29999] = 32'hFFFFFFF1;
    // rom_array[30000] = 32'hFFFFFFF1;
    // rom_array[30001] = 32'hFFFFFFF0;
    // rom_array[30002] = 32'hFFFFFFF0;
    // rom_array[30003] = 32'hFFFFFFF0;
    // rom_array[30004] = 32'hFFFFFFF0;
    // rom_array[30005] = 32'hFFFFFFF1;
    // rom_array[30006] = 32'hFFFFFFF1;
    // rom_array[30007] = 32'hFFFFFFF1;
    // rom_array[30008] = 32'hFFFFFFF1;
    // rom_array[30009] = 32'hFFFFFFF0;
    // rom_array[30010] = 32'hFFFFFFF0;
    // rom_array[30011] = 32'hFFFFFFF1;
    // rom_array[30012] = 32'hFFFFFFF1;
    // rom_array[30013] = 32'hFFFFFFF0;
    // rom_array[30014] = 32'hFFFFFFF0;
    // rom_array[30015] = 32'hFFFFFFF1;
    // rom_array[30016] = 32'hFFFFFFF1;
    // rom_array[30017] = 32'hFFFFFFF0;
    // rom_array[30018] = 32'hFFFFFFF0;
    // rom_array[30019] = 32'hFFFFFFF1;
    // rom_array[30020] = 32'hFFFFFFF1;
    // rom_array[30021] = 32'hFFFFFFF0;
    // rom_array[30022] = 32'hFFFFFFF0;
    // rom_array[30023] = 32'hFFFFFFF1;
    // rom_array[30024] = 32'hFFFFFFF1;
    // rom_array[30025] = 32'hFFFFFFF0;
    // rom_array[30026] = 32'hFFFFFFF0;
    // rom_array[30027] = 32'hFFFFFFF0;
    // rom_array[30028] = 32'hFFFFFFF0;
    // rom_array[30029] = 32'hFFFFFFF1;
    // rom_array[30030] = 32'hFFFFFFF1;
    // rom_array[30031] = 32'hFFFFFFF1;
    // rom_array[30032] = 32'hFFFFFFF1;
    // rom_array[30033] = 32'hFFFFFFF0;
    // rom_array[30034] = 32'hFFFFFFF0;
    // rom_array[30035] = 32'hFFFFFFF0;
    // rom_array[30036] = 32'hFFFFFFF0;
    // rom_array[30037] = 32'hFFFFFFF1;
    // rom_array[30038] = 32'hFFFFFFF1;
    // rom_array[30039] = 32'hFFFFFFF1;
    // rom_array[30040] = 32'hFFFFFFF1;
    // rom_array[30041] = 32'hFFFFFFF0;
    // rom_array[30042] = 32'hFFFFFFF0;
    // rom_array[30043] = 32'hFFFFFFF0;
    // rom_array[30044] = 32'hFFFFFFF0;
    // rom_array[30045] = 32'hFFFFFFF1;
    // rom_array[30046] = 32'hFFFFFFF1;
    // rom_array[30047] = 32'hFFFFFFF1;
    // rom_array[30048] = 32'hFFFFFFF1;
    // rom_array[30049] = 32'hFFFFFFF0;
    // rom_array[30050] = 32'hFFFFFFF0;
    // rom_array[30051] = 32'hFFFFFFF0;
    // rom_array[30052] = 32'hFFFFFFF0;
    // rom_array[30053] = 32'hFFFFFFF1;
    // rom_array[30054] = 32'hFFFFFFF1;
    // rom_array[30055] = 32'hFFFFFFF1;
    // rom_array[30056] = 32'hFFFFFFF1;
    // rom_array[30057] = 32'hFFFFFFF0;
    // rom_array[30058] = 32'hFFFFFFF0;
    // rom_array[30059] = 32'hFFFFFFF1;
    // rom_array[30060] = 32'hFFFFFFF1;
    // rom_array[30061] = 32'hFFFFFFF0;
    // rom_array[30062] = 32'hFFFFFFF0;
    // rom_array[30063] = 32'hFFFFFFF1;
    // rom_array[30064] = 32'hFFFFFFF1;
    // rom_array[30065] = 32'hFFFFFFF0;
    // rom_array[30066] = 32'hFFFFFFF0;
    // rom_array[30067] = 32'hFFFFFFF1;
    // rom_array[30068] = 32'hFFFFFFF1;
    // rom_array[30069] = 32'hFFFFFFF0;
    // rom_array[30070] = 32'hFFFFFFF0;
    // rom_array[30071] = 32'hFFFFFFF1;
    // rom_array[30072] = 32'hFFFFFFF1;
    // rom_array[30073] = 32'hFFFFFFF0;
    // rom_array[30074] = 32'hFFFFFFF0;
    // rom_array[30075] = 32'hFFFFFFF1;
    // rom_array[30076] = 32'hFFFFFFF1;
    // rom_array[30077] = 32'hFFFFFFF0;
    // rom_array[30078] = 32'hFFFFFFF0;
    // rom_array[30079] = 32'hFFFFFFF1;
    // rom_array[30080] = 32'hFFFFFFF1;
    // rom_array[30081] = 32'hFFFFFFF0;
    // rom_array[30082] = 32'hFFFFFFF0;
    // rom_array[30083] = 32'hFFFFFFF1;
    // rom_array[30084] = 32'hFFFFFFF1;
    // rom_array[30085] = 32'hFFFFFFF0;
    // rom_array[30086] = 32'hFFFFFFF0;
    // rom_array[30087] = 32'hFFFFFFF1;
    // rom_array[30088] = 32'hFFFFFFF1;
    // rom_array[30089] = 32'hFFFFFFF0;
    // rom_array[30090] = 32'hFFFFFFF0;
    // rom_array[30091] = 32'hFFFFFFF1;
    // rom_array[30092] = 32'hFFFFFFF1;
    // rom_array[30093] = 32'hFFFFFFF0;
    // rom_array[30094] = 32'hFFFFFFF0;
    // rom_array[30095] = 32'hFFFFFFF0;
    // rom_array[30096] = 32'hFFFFFFF0;
    // rom_array[30097] = 32'hFFFFFFF0;
    // rom_array[30098] = 32'hFFFFFFF0;
    // rom_array[30099] = 32'hFFFFFFF1;
    // rom_array[30100] = 32'hFFFFFFF1;
    // rom_array[30101] = 32'hFFFFFFF0;
    // rom_array[30102] = 32'hFFFFFFF0;
    // rom_array[30103] = 32'hFFFFFFF0;
    // rom_array[30104] = 32'hFFFFFFF0;
    // rom_array[30105] = 32'hFFFFFFF1;
    // rom_array[30106] = 32'hFFFFFFF1;
    // rom_array[30107] = 32'hFFFFFFF1;
    // rom_array[30108] = 32'hFFFFFFF1;
    // rom_array[30109] = 32'hFFFFFFF0;
    // rom_array[30110] = 32'hFFFFFFF0;
    // rom_array[30111] = 32'hFFFFFFF0;
    // rom_array[30112] = 32'hFFFFFFF0;
    // rom_array[30113] = 32'hFFFFFFF1;
    // rom_array[30114] = 32'hFFFFFFF1;
    // rom_array[30115] = 32'hFFFFFFF1;
    // rom_array[30116] = 32'hFFFFFFF1;
    // rom_array[30117] = 32'hFFFFFFF0;
    // rom_array[30118] = 32'hFFFFFFF0;
    // rom_array[30119] = 32'hFFFFFFF0;
    // rom_array[30120] = 32'hFFFFFFF0;
    // rom_array[30121] = 32'hFFFFFFF1;
    // rom_array[30122] = 32'hFFFFFFF1;
    // rom_array[30123] = 32'hFFFFFFF1;
    // rom_array[30124] = 32'hFFFFFFF1;
    // rom_array[30125] = 32'hFFFFFFF0;
    // rom_array[30126] = 32'hFFFFFFF0;
    // rom_array[30127] = 32'hFFFFFFF0;
    // rom_array[30128] = 32'hFFFFFFF0;
    // rom_array[30129] = 32'hFFFFFFF1;
    // rom_array[30130] = 32'hFFFFFFF1;
    // rom_array[30131] = 32'hFFFFFFF1;
    // rom_array[30132] = 32'hFFFFFFF1;
    // rom_array[30133] = 32'hFFFFFFF0;
    // rom_array[30134] = 32'hFFFFFFF0;
    // rom_array[30135] = 32'hFFFFFFF0;
    // rom_array[30136] = 32'hFFFFFFF0;
    // rom_array[30137] = 32'hFFFFFFF1;
    // rom_array[30138] = 32'hFFFFFFF1;
    // rom_array[30139] = 32'hFFFFFFF1;
    // rom_array[30140] = 32'hFFFFFFF1;
    // rom_array[30141] = 32'hFFFFFFF0;
    // rom_array[30142] = 32'hFFFFFFF0;
    // rom_array[30143] = 32'hFFFFFFF0;
    // rom_array[30144] = 32'hFFFFFFF0;
    // rom_array[30145] = 32'hFFFFFFF1;
    // rom_array[30146] = 32'hFFFFFFF1;
    // rom_array[30147] = 32'hFFFFFFF1;
    // rom_array[30148] = 32'hFFFFFFF1;
    // rom_array[30149] = 32'hFFFFFFF0;
    // rom_array[30150] = 32'hFFFFFFF0;
    // rom_array[30151] = 32'hFFFFFFF0;
    // rom_array[30152] = 32'hFFFFFFF0;
    // rom_array[30153] = 32'hFFFFFFF0;
    // rom_array[30154] = 32'hFFFFFFF0;
    // rom_array[30155] = 32'hFFFFFFF0;
    // rom_array[30156] = 32'hFFFFFFF0;
    // rom_array[30157] = 32'hFFFFFFF1;
    // rom_array[30158] = 32'hFFFFFFF1;
    // rom_array[30159] = 32'hFFFFFFF1;
    // rom_array[30160] = 32'hFFFFFFF1;
    // rom_array[30161] = 32'hFFFFFFF0;
    // rom_array[30162] = 32'hFFFFFFF0;
    // rom_array[30163] = 32'hFFFFFFF0;
    // rom_array[30164] = 32'hFFFFFFF0;
    // rom_array[30165] = 32'hFFFFFFF1;
    // rom_array[30166] = 32'hFFFFFFF1;
    // rom_array[30167] = 32'hFFFFFFF1;
    // rom_array[30168] = 32'hFFFFFFF1;
    // rom_array[30169] = 32'hFFFFFFF0;
    // rom_array[30170] = 32'hFFFFFFF0;
    // rom_array[30171] = 32'hFFFFFFF0;
    // rom_array[30172] = 32'hFFFFFFF0;
    // rom_array[30173] = 32'hFFFFFFF1;
    // rom_array[30174] = 32'hFFFFFFF1;
    // rom_array[30175] = 32'hFFFFFFF1;
    // rom_array[30176] = 32'hFFFFFFF1;
    // rom_array[30177] = 32'hFFFFFFF0;
    // rom_array[30178] = 32'hFFFFFFF0;
    // rom_array[30179] = 32'hFFFFFFF0;
    // rom_array[30180] = 32'hFFFFFFF0;
    // rom_array[30181] = 32'hFFFFFFF1;
    // rom_array[30182] = 32'hFFFFFFF1;
    // rom_array[30183] = 32'hFFFFFFF1;
    // rom_array[30184] = 32'hFFFFFFF1;
    // rom_array[30185] = 32'hFFFFFFF0;
    // rom_array[30186] = 32'hFFFFFFF0;
    // rom_array[30187] = 32'hFFFFFFF0;
    // rom_array[30188] = 32'hFFFFFFF0;
    // rom_array[30189] = 32'hFFFFFFF1;
    // rom_array[30190] = 32'hFFFFFFF1;
    // rom_array[30191] = 32'hFFFFFFF1;
    // rom_array[30192] = 32'hFFFFFFF1;
    // rom_array[30193] = 32'hFFFFFFF0;
    // rom_array[30194] = 32'hFFFFFFF0;
    // rom_array[30195] = 32'hFFFFFFF0;
    // rom_array[30196] = 32'hFFFFFFF0;
    // rom_array[30197] = 32'hFFFFFFF1;
    // rom_array[30198] = 32'hFFFFFFF1;
    // rom_array[30199] = 32'hFFFFFFF1;
    // rom_array[30200] = 32'hFFFFFFF1;
    // rom_array[30201] = 32'hFFFFFFF0;
    // rom_array[30202] = 32'hFFFFFFF0;
    // rom_array[30203] = 32'hFFFFFFF0;
    // rom_array[30204] = 32'hFFFFFFF0;
    // rom_array[30205] = 32'hFFFFFFF1;
    // rom_array[30206] = 32'hFFFFFFF1;
    // rom_array[30207] = 32'hFFFFFFF1;
    // rom_array[30208] = 32'hFFFFFFF1;
    // rom_array[30209] = 32'hFFFFFFF0;
    // rom_array[30210] = 32'hFFFFFFF0;
    // rom_array[30211] = 32'hFFFFFFF0;
    // rom_array[30212] = 32'hFFFFFFF0;
    // rom_array[30213] = 32'hFFFFFFF1;
    // rom_array[30214] = 32'hFFFFFFF1;
    // rom_array[30215] = 32'hFFFFFFF1;
    // rom_array[30216] = 32'hFFFFFFF1;
    // rom_array[30217] = 32'hFFFFFFF0;
    // rom_array[30218] = 32'hFFFFFFF0;
    // rom_array[30219] = 32'hFFFFFFF0;
    // rom_array[30220] = 32'hFFFFFFF0;
    // rom_array[30221] = 32'hFFFFFFF1;
    // rom_array[30222] = 32'hFFFFFFF1;
    // rom_array[30223] = 32'hFFFFFFF1;
    // rom_array[30224] = 32'hFFFFFFF1;
    // rom_array[30225] = 32'hFFFFFFF0;
    // rom_array[30226] = 32'hFFFFFFF0;
    // rom_array[30227] = 32'hFFFFFFF0;
    // rom_array[30228] = 32'hFFFFFFF0;
    // rom_array[30229] = 32'hFFFFFFF1;
    // rom_array[30230] = 32'hFFFFFFF1;
    // rom_array[30231] = 32'hFFFFFFF1;
    // rom_array[30232] = 32'hFFFFFFF1;
    // rom_array[30233] = 32'hFFFFFFF0;
    // rom_array[30234] = 32'hFFFFFFF0;
    // rom_array[30235] = 32'hFFFFFFF0;
    // rom_array[30236] = 32'hFFFFFFF0;
    // rom_array[30237] = 32'hFFFFFFF1;
    // rom_array[30238] = 32'hFFFFFFF1;
    // rom_array[30239] = 32'hFFFFFFF1;
    // rom_array[30240] = 32'hFFFFFFF1;
    // rom_array[30241] = 32'hFFFFFFF0;
    // rom_array[30242] = 32'hFFFFFFF0;
    // rom_array[30243] = 32'hFFFFFFF0;
    // rom_array[30244] = 32'hFFFFFFF0;
    // rom_array[30245] = 32'hFFFFFFF1;
    // rom_array[30246] = 32'hFFFFFFF1;
    // rom_array[30247] = 32'hFFFFFFF1;
    // rom_array[30248] = 32'hFFFFFFF1;
    // rom_array[30249] = 32'hFFFFFFF0;
    // rom_array[30250] = 32'hFFFFFFF0;
    // rom_array[30251] = 32'hFFFFFFF0;
    // rom_array[30252] = 32'hFFFFFFF0;
    // rom_array[30253] = 32'hFFFFFFF1;
    // rom_array[30254] = 32'hFFFFFFF1;
    // rom_array[30255] = 32'hFFFFFFF1;
    // rom_array[30256] = 32'hFFFFFFF1;
    // rom_array[30257] = 32'hFFFFFFF0;
    // rom_array[30258] = 32'hFFFFFFF0;
    // rom_array[30259] = 32'hFFFFFFF0;
    // rom_array[30260] = 32'hFFFFFFF0;
    // rom_array[30261] = 32'hFFFFFFF1;
    // rom_array[30262] = 32'hFFFFFFF1;
    // rom_array[30263] = 32'hFFFFFFF1;
    // rom_array[30264] = 32'hFFFFFFF1;
    // rom_array[30265] = 32'hFFFFFFF0;
    // rom_array[30266] = 32'hFFFFFFF0;
    // rom_array[30267] = 32'hFFFFFFF0;
    // rom_array[30268] = 32'hFFFFFFF0;
    // rom_array[30269] = 32'hFFFFFFF1;
    // rom_array[30270] = 32'hFFFFFFF1;
    // rom_array[30271] = 32'hFFFFFFF1;
    // rom_array[30272] = 32'hFFFFFFF1;
    // rom_array[30273] = 32'hFFFFFFF0;
    // rom_array[30274] = 32'hFFFFFFF0;
    // rom_array[30275] = 32'hFFFFFFF0;
    // rom_array[30276] = 32'hFFFFFFF0;
    // rom_array[30277] = 32'hFFFFFFF1;
    // rom_array[30278] = 32'hFFFFFFF1;
    // rom_array[30279] = 32'hFFFFFFF1;
    // rom_array[30280] = 32'hFFFFFFF1;
    // rom_array[30281] = 32'hFFFFFFF1;
    // rom_array[30282] = 32'hFFFFFFF1;
    // rom_array[30283] = 32'hFFFFFFF1;
    // rom_array[30284] = 32'hFFFFFFF1;
    // rom_array[30285] = 32'hFFFFFFF0;
    // rom_array[30286] = 32'hFFFFFFF0;
    // rom_array[30287] = 32'hFFFFFFF0;
    // rom_array[30288] = 32'hFFFFFFF0;
    // rom_array[30289] = 32'hFFFFFFF1;
    // rom_array[30290] = 32'hFFFFFFF1;
    // rom_array[30291] = 32'hFFFFFFF1;
    // rom_array[30292] = 32'hFFFFFFF1;
    // rom_array[30293] = 32'hFFFFFFF0;
    // rom_array[30294] = 32'hFFFFFFF0;
    // rom_array[30295] = 32'hFFFFFFF0;
    // rom_array[30296] = 32'hFFFFFFF0;
    // rom_array[30297] = 32'hFFFFFFF1;
    // rom_array[30298] = 32'hFFFFFFF1;
    // rom_array[30299] = 32'hFFFFFFF1;
    // rom_array[30300] = 32'hFFFFFFF1;
    // rom_array[30301] = 32'hFFFFFFF0;
    // rom_array[30302] = 32'hFFFFFFF0;
    // rom_array[30303] = 32'hFFFFFFF0;
    // rom_array[30304] = 32'hFFFFFFF0;
    // rom_array[30305] = 32'hFFFFFFF1;
    // rom_array[30306] = 32'hFFFFFFF1;
    // rom_array[30307] = 32'hFFFFFFF1;
    // rom_array[30308] = 32'hFFFFFFF1;
    // rom_array[30309] = 32'hFFFFFFF0;
    // rom_array[30310] = 32'hFFFFFFF0;
    // rom_array[30311] = 32'hFFFFFFF0;
    // rom_array[30312] = 32'hFFFFFFF0;
    // rom_array[30313] = 32'hFFFFFFF1;
    // rom_array[30314] = 32'hFFFFFFF1;
    // rom_array[30315] = 32'hFFFFFFF1;
    // rom_array[30316] = 32'hFFFFFFF1;
    // rom_array[30317] = 32'hFFFFFFF0;
    // rom_array[30318] = 32'hFFFFFFF0;
    // rom_array[30319] = 32'hFFFFFFF0;
    // rom_array[30320] = 32'hFFFFFFF0;
    // rom_array[30321] = 32'hFFFFFFF1;
    // rom_array[30322] = 32'hFFFFFFF1;
    // rom_array[30323] = 32'hFFFFFFF1;
    // rom_array[30324] = 32'hFFFFFFF1;
    // rom_array[30325] = 32'hFFFFFFF0;
    // rom_array[30326] = 32'hFFFFFFF0;
    // rom_array[30327] = 32'hFFFFFFF0;
    // rom_array[30328] = 32'hFFFFFFF0;
    // rom_array[30329] = 32'hFFFFFFF1;
    // rom_array[30330] = 32'hFFFFFFF1;
    // rom_array[30331] = 32'hFFFFFFF1;
    // rom_array[30332] = 32'hFFFFFFF1;
    // rom_array[30333] = 32'hFFFFFFF0;
    // rom_array[30334] = 32'hFFFFFFF0;
    // rom_array[30335] = 32'hFFFFFFF0;
    // rom_array[30336] = 32'hFFFFFFF0;
    // rom_array[30337] = 32'hFFFFFFF1;
    // rom_array[30338] = 32'hFFFFFFF1;
    // rom_array[30339] = 32'hFFFFFFF1;
    // rom_array[30340] = 32'hFFFFFFF1;
    // rom_array[30341] = 32'hFFFFFFF0;
    // rom_array[30342] = 32'hFFFFFFF0;
    // rom_array[30343] = 32'hFFFFFFF0;
    // rom_array[30344] = 32'hFFFFFFF0;
    // rom_array[30345] = 32'hFFFFFFF1;
    // rom_array[30346] = 32'hFFFFFFF1;
    // rom_array[30347] = 32'hFFFFFFF1;
    // rom_array[30348] = 32'hFFFFFFF1;
    // rom_array[30349] = 32'hFFFFFFF0;
    // rom_array[30350] = 32'hFFFFFFF0;
    // rom_array[30351] = 32'hFFFFFFF1;
    // rom_array[30352] = 32'hFFFFFFF1;
    // rom_array[30353] = 32'hFFFFFFF1;
    // rom_array[30354] = 32'hFFFFFFF1;
    // rom_array[30355] = 32'hFFFFFFF1;
    // rom_array[30356] = 32'hFFFFFFF1;
    // rom_array[30357] = 32'hFFFFFFF0;
    // rom_array[30358] = 32'hFFFFFFF0;
    // rom_array[30359] = 32'hFFFFFFF1;
    // rom_array[30360] = 32'hFFFFFFF1;
    // rom_array[30361] = 32'hFFFFFFF1;
    // rom_array[30362] = 32'hFFFFFFF1;
    // rom_array[30363] = 32'hFFFFFFF1;
    // rom_array[30364] = 32'hFFFFFFF1;
    // rom_array[30365] = 32'hFFFFFFF1;
    // rom_array[30366] = 32'hFFFFFFF1;
    // rom_array[30367] = 32'hFFFFFFF1;
    // rom_array[30368] = 32'hFFFFFFF1;
    // rom_array[30369] = 32'hFFFFFFF1;
    // rom_array[30370] = 32'hFFFFFFF1;
    // rom_array[30371] = 32'hFFFFFFF1;
    // rom_array[30372] = 32'hFFFFFFF1;
    // rom_array[30373] = 32'hFFFFFFF1;
    // rom_array[30374] = 32'hFFFFFFF1;
    // rom_array[30375] = 32'hFFFFFFF1;
    // rom_array[30376] = 32'hFFFFFFF1;
    // rom_array[30377] = 32'hFFFFFFF0;
    // rom_array[30378] = 32'hFFFFFFF0;
    // rom_array[30379] = 32'hFFFFFFF1;
    // rom_array[30380] = 32'hFFFFFFF1;
    // rom_array[30381] = 32'hFFFFFFF0;
    // rom_array[30382] = 32'hFFFFFFF0;
    // rom_array[30383] = 32'hFFFFFFF1;
    // rom_array[30384] = 32'hFFFFFFF1;
    // rom_array[30385] = 32'hFFFFFFF0;
    // rom_array[30386] = 32'hFFFFFFF0;
    // rom_array[30387] = 32'hFFFFFFF1;
    // rom_array[30388] = 32'hFFFFFFF1;
    // rom_array[30389] = 32'hFFFFFFF0;
    // rom_array[30390] = 32'hFFFFFFF0;
    // rom_array[30391] = 32'hFFFFFFF1;
    // rom_array[30392] = 32'hFFFFFFF1;
    // rom_array[30393] = 32'hFFFFFFF1;
    // rom_array[30394] = 32'hFFFFFFF1;
    // rom_array[30395] = 32'hFFFFFFF1;
    // rom_array[30396] = 32'hFFFFFFF1;
    // rom_array[30397] = 32'hFFFFFFF1;
    // rom_array[30398] = 32'hFFFFFFF1;
    // rom_array[30399] = 32'hFFFFFFF1;
    // rom_array[30400] = 32'hFFFFFFF1;
    // rom_array[30401] = 32'hFFFFFFF1;
    // rom_array[30402] = 32'hFFFFFFF1;
    // rom_array[30403] = 32'hFFFFFFF1;
    // rom_array[30404] = 32'hFFFFFFF1;
    // rom_array[30405] = 32'hFFFFFFF1;
    // rom_array[30406] = 32'hFFFFFFF1;
    // rom_array[30407] = 32'hFFFFFFF1;
    // rom_array[30408] = 32'hFFFFFFF1;
    // rom_array[30409] = 32'hFFFFFFF1;
    // rom_array[30410] = 32'hFFFFFFF1;
    // rom_array[30411] = 32'hFFFFFFF1;
    // rom_array[30412] = 32'hFFFFFFF1;
    // rom_array[30413] = 32'hFFFFFFF1;
    // rom_array[30414] = 32'hFFFFFFF1;
    // rom_array[30415] = 32'hFFFFFFF1;
    // rom_array[30416] = 32'hFFFFFFF1;
    // rom_array[30417] = 32'hFFFFFFF1;
    // rom_array[30418] = 32'hFFFFFFF1;
    // rom_array[30419] = 32'hFFFFFFF1;
    // rom_array[30420] = 32'hFFFFFFF1;
    // rom_array[30421] = 32'hFFFFFFF1;
    // rom_array[30422] = 32'hFFFFFFF1;
    // rom_array[30423] = 32'hFFFFFFF1;
    // rom_array[30424] = 32'hFFFFFFF1;
    // rom_array[30425] = 32'hFFFFFFF0;
    // rom_array[30426] = 32'hFFFFFFF0;
    // rom_array[30427] = 32'hFFFFFFF1;
    // rom_array[30428] = 32'hFFFFFFF1;
    // rom_array[30429] = 32'hFFFFFFF0;
    // rom_array[30430] = 32'hFFFFFFF0;
    // rom_array[30431] = 32'hFFFFFFF1;
    // rom_array[30432] = 32'hFFFFFFF1;
    // rom_array[30433] = 32'hFFFFFFF0;
    // rom_array[30434] = 32'hFFFFFFF0;
    // rom_array[30435] = 32'hFFFFFFF1;
    // rom_array[30436] = 32'hFFFFFFF1;
    // rom_array[30437] = 32'hFFFFFFF0;
    // rom_array[30438] = 32'hFFFFFFF0;
    // rom_array[30439] = 32'hFFFFFFF1;
    // rom_array[30440] = 32'hFFFFFFF1;
    // rom_array[30441] = 32'hFFFFFFF1;
    // rom_array[30442] = 32'hFFFFFFF1;
    // rom_array[30443] = 32'hFFFFFFF1;
    // rom_array[30444] = 32'hFFFFFFF1;
    // rom_array[30445] = 32'hFFFFFFF1;
    // rom_array[30446] = 32'hFFFFFFF1;
    // rom_array[30447] = 32'hFFFFFFF1;
    // rom_array[30448] = 32'hFFFFFFF1;
    // rom_array[30449] = 32'hFFFFFFF1;
    // rom_array[30450] = 32'hFFFFFFF1;
    // rom_array[30451] = 32'hFFFFFFF1;
    // rom_array[30452] = 32'hFFFFFFF1;
    // rom_array[30453] = 32'hFFFFFFF1;
    // rom_array[30454] = 32'hFFFFFFF1;
    // rom_array[30455] = 32'hFFFFFFF1;
    // rom_array[30456] = 32'hFFFFFFF1;
    // rom_array[30457] = 32'hFFFFFFF0;
    // rom_array[30458] = 32'hFFFFFFF0;
    // rom_array[30459] = 32'hFFFFFFF1;
    // rom_array[30460] = 32'hFFFFFFF1;
    // rom_array[30461] = 32'hFFFFFFF0;
    // rom_array[30462] = 32'hFFFFFFF0;
    // rom_array[30463] = 32'hFFFFFFF1;
    // rom_array[30464] = 32'hFFFFFFF1;
    // rom_array[30465] = 32'hFFFFFFF0;
    // rom_array[30466] = 32'hFFFFFFF0;
    // rom_array[30467] = 32'hFFFFFFF1;
    // rom_array[30468] = 32'hFFFFFFF1;
    // rom_array[30469] = 32'hFFFFFFF0;
    // rom_array[30470] = 32'hFFFFFFF0;
    // rom_array[30471] = 32'hFFFFFFF1;
    // rom_array[30472] = 32'hFFFFFFF1;
    // rom_array[30473] = 32'hFFFFFFF1;
    // rom_array[30474] = 32'hFFFFFFF1;
    // rom_array[30475] = 32'hFFFFFFF1;
    // rom_array[30476] = 32'hFFFFFFF1;
    // rom_array[30477] = 32'hFFFFFFF1;
    // rom_array[30478] = 32'hFFFFFFF1;
    // rom_array[30479] = 32'hFFFFFFF1;
    // rom_array[30480] = 32'hFFFFFFF1;
    // rom_array[30481] = 32'hFFFFFFF1;
    // rom_array[30482] = 32'hFFFFFFF1;
    // rom_array[30483] = 32'hFFFFFFF1;
    // rom_array[30484] = 32'hFFFFFFF1;
    // rom_array[30485] = 32'hFFFFFFF1;
    // rom_array[30486] = 32'hFFFFFFF1;
    // rom_array[30487] = 32'hFFFFFFF1;
    // rom_array[30488] = 32'hFFFFFFF1;
    // rom_array[30489] = 32'hFFFFFFF1;
    // rom_array[30490] = 32'hFFFFFFF1;
    // rom_array[30491] = 32'hFFFFFFF1;
    // rom_array[30492] = 32'hFFFFFFF1;
    // rom_array[30493] = 32'hFFFFFFF1;
    // rom_array[30494] = 32'hFFFFFFF1;
    // rom_array[30495] = 32'hFFFFFFF1;
    // rom_array[30496] = 32'hFFFFFFF1;
    // rom_array[30497] = 32'hFFFFFFF1;
    // rom_array[30498] = 32'hFFFFFFF1;
    // rom_array[30499] = 32'hFFFFFFF1;
    // rom_array[30500] = 32'hFFFFFFF1;
    // rom_array[30501] = 32'hFFFFFFF1;
    // rom_array[30502] = 32'hFFFFFFF1;
    // rom_array[30503] = 32'hFFFFFFF1;
    // rom_array[30504] = 32'hFFFFFFF1;
    // rom_array[30505] = 32'hFFFFFFF1;
    // rom_array[30506] = 32'hFFFFFFF1;
    // rom_array[30507] = 32'hFFFFFFF1;
    // rom_array[30508] = 32'hFFFFFFF1;
    // rom_array[30509] = 32'hFFFFFFF1;
    // rom_array[30510] = 32'hFFFFFFF1;
    // rom_array[30511] = 32'hFFFFFFF1;
    // rom_array[30512] = 32'hFFFFFFF1;
    // rom_array[30513] = 32'hFFFFFFF1;
    // rom_array[30514] = 32'hFFFFFFF1;
    // rom_array[30515] = 32'hFFFFFFF1;
    // rom_array[30516] = 32'hFFFFFFF1;
    // rom_array[30517] = 32'hFFFFFFF1;
    // rom_array[30518] = 32'hFFFFFFF1;
    // rom_array[30519] = 32'hFFFFFFF1;
    // rom_array[30520] = 32'hFFFFFFF1;
    // rom_array[30521] = 32'hFFFFFFF0;
    // rom_array[30522] = 32'hFFFFFFF0;
    // rom_array[30523] = 32'hFFFFFFF1;
    // rom_array[30524] = 32'hFFFFFFF1;
    // rom_array[30525] = 32'hFFFFFFF0;
    // rom_array[30526] = 32'hFFFFFFF0;
    // rom_array[30527] = 32'hFFFFFFF1;
    // rom_array[30528] = 32'hFFFFFFF1;
    // rom_array[30529] = 32'hFFFFFFF0;
    // rom_array[30530] = 32'hFFFFFFF0;
    // rom_array[30531] = 32'hFFFFFFF1;
    // rom_array[30532] = 32'hFFFFFFF1;
    // rom_array[30533] = 32'hFFFFFFF0;
    // rom_array[30534] = 32'hFFFFFFF0;
    // rom_array[30535] = 32'hFFFFFFF1;
    // rom_array[30536] = 32'hFFFFFFF1;
    // rom_array[30537] = 32'hFFFFFFF1;
    // rom_array[30538] = 32'hFFFFFFF1;
    // rom_array[30539] = 32'hFFFFFFF1;
    // rom_array[30540] = 32'hFFFFFFF1;
    // rom_array[30541] = 32'hFFFFFFF1;
    // rom_array[30542] = 32'hFFFFFFF1;
    // rom_array[30543] = 32'hFFFFFFF1;
    // rom_array[30544] = 32'hFFFFFFF1;
    // rom_array[30545] = 32'hFFFFFFF1;
    // rom_array[30546] = 32'hFFFFFFF1;
    // rom_array[30547] = 32'hFFFFFFF1;
    // rom_array[30548] = 32'hFFFFFFF1;
    // rom_array[30549] = 32'hFFFFFFF1;
    // rom_array[30550] = 32'hFFFFFFF1;
    // rom_array[30551] = 32'hFFFFFFF1;
    // rom_array[30552] = 32'hFFFFFFF1;
    // rom_array[30553] = 32'hFFFFFFF0;
    // rom_array[30554] = 32'hFFFFFFF0;
    // rom_array[30555] = 32'hFFFFFFF1;
    // rom_array[30556] = 32'hFFFFFFF1;
    // rom_array[30557] = 32'hFFFFFFF0;
    // rom_array[30558] = 32'hFFFFFFF0;
    // rom_array[30559] = 32'hFFFFFFF1;
    // rom_array[30560] = 32'hFFFFFFF1;
    // rom_array[30561] = 32'hFFFFFFF0;
    // rom_array[30562] = 32'hFFFFFFF0;
    // rom_array[30563] = 32'hFFFFFFF1;
    // rom_array[30564] = 32'hFFFFFFF1;
    // rom_array[30565] = 32'hFFFFFFF0;
    // rom_array[30566] = 32'hFFFFFFF0;
    // rom_array[30567] = 32'hFFFFFFF1;
    // rom_array[30568] = 32'hFFFFFFF1;
    // rom_array[30569] = 32'hFFFFFFF1;
    // rom_array[30570] = 32'hFFFFFFF1;
    // rom_array[30571] = 32'hFFFFFFF1;
    // rom_array[30572] = 32'hFFFFFFF1;
    // rom_array[30573] = 32'hFFFFFFF1;
    // rom_array[30574] = 32'hFFFFFFF1;
    // rom_array[30575] = 32'hFFFFFFF1;
    // rom_array[30576] = 32'hFFFFFFF1;
    // rom_array[30577] = 32'hFFFFFFF1;
    // rom_array[30578] = 32'hFFFFFFF1;
    // rom_array[30579] = 32'hFFFFFFF1;
    // rom_array[30580] = 32'hFFFFFFF1;
    // rom_array[30581] = 32'hFFFFFFF1;
    // rom_array[30582] = 32'hFFFFFFF1;
    // rom_array[30583] = 32'hFFFFFFF1;
    // rom_array[30584] = 32'hFFFFFFF1;
    // rom_array[30585] = 32'hFFFFFFF0;
    // rom_array[30586] = 32'hFFFFFFF0;
    // rom_array[30587] = 32'hFFFFFFF0;
    // rom_array[30588] = 32'hFFFFFFF0;
    // rom_array[30589] = 32'hFFFFFFF1;
    // rom_array[30590] = 32'hFFFFFFF1;
    // rom_array[30591] = 32'hFFFFFFF1;
    // rom_array[30592] = 32'hFFFFFFF1;
    // rom_array[30593] = 32'hFFFFFFF0;
    // rom_array[30594] = 32'hFFFFFFF0;
    // rom_array[30595] = 32'hFFFFFFF0;
    // rom_array[30596] = 32'hFFFFFFF0;
    // rom_array[30597] = 32'hFFFFFFF1;
    // rom_array[30598] = 32'hFFFFFFF1;
    // rom_array[30599] = 32'hFFFFFFF1;
    // rom_array[30600] = 32'hFFFFFFF1;
    // rom_array[30601] = 32'hFFFFFFF0;
    // rom_array[30602] = 32'hFFFFFFF0;
    // rom_array[30603] = 32'hFFFFFFF1;
    // rom_array[30604] = 32'hFFFFFFF1;
    // rom_array[30605] = 32'hFFFFFFF0;
    // rom_array[30606] = 32'hFFFFFFF0;
    // rom_array[30607] = 32'hFFFFFFF1;
    // rom_array[30608] = 32'hFFFFFFF1;
    // rom_array[30609] = 32'hFFFFFFF0;
    // rom_array[30610] = 32'hFFFFFFF0;
    // rom_array[30611] = 32'hFFFFFFF1;
    // rom_array[30612] = 32'hFFFFFFF1;
    // rom_array[30613] = 32'hFFFFFFF0;
    // rom_array[30614] = 32'hFFFFFFF0;
    // rom_array[30615] = 32'hFFFFFFF1;
    // rom_array[30616] = 32'hFFFFFFF1;
    // rom_array[30617] = 32'hFFFFFFF1;
    // rom_array[30618] = 32'hFFFFFFF1;
    // rom_array[30619] = 32'hFFFFFFF1;
    // rom_array[30620] = 32'hFFFFFFF1;
    // rom_array[30621] = 32'hFFFFFFF1;
    // rom_array[30622] = 32'hFFFFFFF1;
    // rom_array[30623] = 32'hFFFFFFF1;
    // rom_array[30624] = 32'hFFFFFFF1;
    // rom_array[30625] = 32'hFFFFFFF1;
    // rom_array[30626] = 32'hFFFFFFF1;
    // rom_array[30627] = 32'hFFFFFFF1;
    // rom_array[30628] = 32'hFFFFFFF1;
    // rom_array[30629] = 32'hFFFFFFF1;
    // rom_array[30630] = 32'hFFFFFFF1;
    // rom_array[30631] = 32'hFFFFFFF1;
    // rom_array[30632] = 32'hFFFFFFF1;
    // rom_array[30633] = 32'hFFFFFFF0;
    // rom_array[30634] = 32'hFFFFFFF0;
    // rom_array[30635] = 32'hFFFFFFF1;
    // rom_array[30636] = 32'hFFFFFFF1;
    // rom_array[30637] = 32'hFFFFFFF0;
    // rom_array[30638] = 32'hFFFFFFF0;
    // rom_array[30639] = 32'hFFFFFFF1;
    // rom_array[30640] = 32'hFFFFFFF1;
    // rom_array[30641] = 32'hFFFFFFF0;
    // rom_array[30642] = 32'hFFFFFFF0;
    // rom_array[30643] = 32'hFFFFFFF1;
    // rom_array[30644] = 32'hFFFFFFF1;
    // rom_array[30645] = 32'hFFFFFFF0;
    // rom_array[30646] = 32'hFFFFFFF0;
    // rom_array[30647] = 32'hFFFFFFF1;
    // rom_array[30648] = 32'hFFFFFFF1;
    // rom_array[30649] = 32'hFFFFFFF1;
    // rom_array[30650] = 32'hFFFFFFF1;
    // rom_array[30651] = 32'hFFFFFFF1;
    // rom_array[30652] = 32'hFFFFFFF1;
    // rom_array[30653] = 32'hFFFFFFF1;
    // rom_array[30654] = 32'hFFFFFFF1;
    // rom_array[30655] = 32'hFFFFFFF1;
    // rom_array[30656] = 32'hFFFFFFF1;
    // rom_array[30657] = 32'hFFFFFFF1;
    // rom_array[30658] = 32'hFFFFFFF1;
    // rom_array[30659] = 32'hFFFFFFF1;
    // rom_array[30660] = 32'hFFFFFFF1;
    // rom_array[30661] = 32'hFFFFFFF1;
    // rom_array[30662] = 32'hFFFFFFF1;
    // rom_array[30663] = 32'hFFFFFFF1;
    // rom_array[30664] = 32'hFFFFFFF1;
    // rom_array[30665] = 32'hFFFFFFF1;
    // rom_array[30666] = 32'hFFFFFFF1;
    // rom_array[30667] = 32'hFFFFFFF1;
    // rom_array[30668] = 32'hFFFFFFF1;
    // rom_array[30669] = 32'hFFFFFFF1;
    // rom_array[30670] = 32'hFFFFFFF1;
    // rom_array[30671] = 32'hFFFFFFF1;
    // rom_array[30672] = 32'hFFFFFFF1;
    // rom_array[30673] = 32'hFFFFFFF1;
    // rom_array[30674] = 32'hFFFFFFF1;
    // rom_array[30675] = 32'hFFFFFFF1;
    // rom_array[30676] = 32'hFFFFFFF1;
    // rom_array[30677] = 32'hFFFFFFF1;
    // rom_array[30678] = 32'hFFFFFFF1;
    // rom_array[30679] = 32'hFFFFFFF1;
    // rom_array[30680] = 32'hFFFFFFF1;
    // rom_array[30681] = 32'hFFFFFFF1;
    // rom_array[30682] = 32'hFFFFFFF1;
    // rom_array[30683] = 32'hFFFFFFF1;
    // rom_array[30684] = 32'hFFFFFFF1;
    // rom_array[30685] = 32'hFFFFFFF1;
    // rom_array[30686] = 32'hFFFFFFF1;
    // rom_array[30687] = 32'hFFFFFFF1;
    // rom_array[30688] = 32'hFFFFFFF1;
    // rom_array[30689] = 32'hFFFFFFF1;
    // rom_array[30690] = 32'hFFFFFFF1;
    // rom_array[30691] = 32'hFFFFFFF1;
    // rom_array[30692] = 32'hFFFFFFF1;
    // rom_array[30693] = 32'hFFFFFFF1;
    // rom_array[30694] = 32'hFFFFFFF1;
    // rom_array[30695] = 32'hFFFFFFF1;
    // rom_array[30696] = 32'hFFFFFFF1;
    // rom_array[30697] = 32'hFFFFFFF1;
    // rom_array[30698] = 32'hFFFFFFF1;
    // rom_array[30699] = 32'hFFFFFFF1;
    // rom_array[30700] = 32'hFFFFFFF1;
    // rom_array[30701] = 32'hFFFFFFF1;
    // rom_array[30702] = 32'hFFFFFFF1;
    // rom_array[30703] = 32'hFFFFFFF1;
    // rom_array[30704] = 32'hFFFFFFF1;
    // rom_array[30705] = 32'hFFFFFFF1;
    // rom_array[30706] = 32'hFFFFFFF1;
    // rom_array[30707] = 32'hFFFFFFF1;
    // rom_array[30708] = 32'hFFFFFFF1;
    // rom_array[30709] = 32'hFFFFFFF1;
    // rom_array[30710] = 32'hFFFFFFF1;
    // rom_array[30711] = 32'hFFFFFFF1;
    // rom_array[30712] = 32'hFFFFFFF1;
    // rom_array[30713] = 32'hFFFFFFF1;
    // rom_array[30714] = 32'hFFFFFFF1;
    // rom_array[30715] = 32'hFFFFFFF1;
    // rom_array[30716] = 32'hFFFFFFF1;
    // rom_array[30717] = 32'hFFFFFFF1;
    // rom_array[30718] = 32'hFFFFFFF1;
    // rom_array[30719] = 32'hFFFFFFF1;
    // rom_array[30720] = 32'hFFFFFFF1;
    // rom_array[30721] = 32'hFFFFFFF1;
    // rom_array[30722] = 32'hFFFFFFF1;
    // rom_array[30723] = 32'hFFFFFFF1;
    // rom_array[30724] = 32'hFFFFFFF1;
    // rom_array[30725] = 32'hFFFFFFF1;
    // rom_array[30726] = 32'hFFFFFFF1;
    // rom_array[30727] = 32'hFFFFFFF1;
    // rom_array[30728] = 32'hFFFFFFF1;
    // rom_array[30729] = 32'hFFFFFFF1;
    // rom_array[30730] = 32'hFFFFFFF1;
    // rom_array[30731] = 32'hFFFFFFF1;
    // rom_array[30732] = 32'hFFFFFFF1;
    // rom_array[30733] = 32'hFFFFFFF1;
    // rom_array[30734] = 32'hFFFFFFF1;
    // rom_array[30735] = 32'hFFFFFFF1;
    // rom_array[30736] = 32'hFFFFFFF1;
    // rom_array[30737] = 32'hFFFFFFF1;
    // rom_array[30738] = 32'hFFFFFFF1;
    // rom_array[30739] = 32'hFFFFFFF1;
    // rom_array[30740] = 32'hFFFFFFF1;
    // rom_array[30741] = 32'hFFFFFFF1;
    // rom_array[30742] = 32'hFFFFFFF1;
    // rom_array[30743] = 32'hFFFFFFF1;
    // rom_array[30744] = 32'hFFFFFFF1;
    // rom_array[30745] = 32'hFFFFFFF1;
    // rom_array[30746] = 32'hFFFFFFF1;
    // rom_array[30747] = 32'hFFFFFFF1;
    // rom_array[30748] = 32'hFFFFFFF1;
    // rom_array[30749] = 32'hFFFFFFF1;
    // rom_array[30750] = 32'hFFFFFFF1;
    // rom_array[30751] = 32'hFFFFFFF1;
    // rom_array[30752] = 32'hFFFFFFF1;
    // rom_array[30753] = 32'hFFFFFFF1;
    // rom_array[30754] = 32'hFFFFFFF1;
    // rom_array[30755] = 32'hFFFFFFF1;
    // rom_array[30756] = 32'hFFFFFFF1;
    // rom_array[30757] = 32'hFFFFFFF1;
    // rom_array[30758] = 32'hFFFFFFF1;
    // rom_array[30759] = 32'hFFFFFFF1;
    // rom_array[30760] = 32'hFFFFFFF1;
    // rom_array[30761] = 32'hFFFFFFF0;
    // rom_array[30762] = 32'hFFFFFFF0;
    // rom_array[30763] = 32'hFFFFFFF1;
    // rom_array[30764] = 32'hFFFFFFF1;
    // rom_array[30765] = 32'hFFFFFFF0;
    // rom_array[30766] = 32'hFFFFFFF0;
    // rom_array[30767] = 32'hFFFFFFF1;
    // rom_array[30768] = 32'hFFFFFFF1;
    // rom_array[30769] = 32'hFFFFFFF0;
    // rom_array[30770] = 32'hFFFFFFF0;
    // rom_array[30771] = 32'hFFFFFFF1;
    // rom_array[30772] = 32'hFFFFFFF1;
    // rom_array[30773] = 32'hFFFFFFF0;
    // rom_array[30774] = 32'hFFFFFFF0;
    // rom_array[30775] = 32'hFFFFFFF1;
    // rom_array[30776] = 32'hFFFFFFF1;
    // rom_array[30777] = 32'hFFFFFFF0;
    // rom_array[30778] = 32'hFFFFFFF0;
    // rom_array[30779] = 32'hFFFFFFF1;
    // rom_array[30780] = 32'hFFFFFFF1;
    // rom_array[30781] = 32'hFFFFFFF0;
    // rom_array[30782] = 32'hFFFFFFF0;
    // rom_array[30783] = 32'hFFFFFFF1;
    // rom_array[30784] = 32'hFFFFFFF1;
    // rom_array[30785] = 32'hFFFFFFF0;
    // rom_array[30786] = 32'hFFFFFFF0;
    // rom_array[30787] = 32'hFFFFFFF1;
    // rom_array[30788] = 32'hFFFFFFF1;
    // rom_array[30789] = 32'hFFFFFFF0;
    // rom_array[30790] = 32'hFFFFFFF0;
    // rom_array[30791] = 32'hFFFFFFF1;
    // rom_array[30792] = 32'hFFFFFFF1;
    // rom_array[30793] = 32'hFFFFFFF1;
    // rom_array[30794] = 32'hFFFFFFF1;
    // rom_array[30795] = 32'hFFFFFFF1;
    // rom_array[30796] = 32'hFFFFFFF1;
    // rom_array[30797] = 32'hFFFFFFF1;
    // rom_array[30798] = 32'hFFFFFFF1;
    // rom_array[30799] = 32'hFFFFFFF1;
    // rom_array[30800] = 32'hFFFFFFF1;
    // rom_array[30801] = 32'hFFFFFFF1;
    // rom_array[30802] = 32'hFFFFFFF1;
    // rom_array[30803] = 32'hFFFFFFF1;
    // rom_array[30804] = 32'hFFFFFFF1;
    // rom_array[30805] = 32'hFFFFFFF1;
    // rom_array[30806] = 32'hFFFFFFF1;
    // rom_array[30807] = 32'hFFFFFFF1;
    // rom_array[30808] = 32'hFFFFFFF1;
    // rom_array[30809] = 32'hFFFFFFF1;
    // rom_array[30810] = 32'hFFFFFFF1;
    // rom_array[30811] = 32'hFFFFFFF1;
    // rom_array[30812] = 32'hFFFFFFF1;
    // rom_array[30813] = 32'hFFFFFFF1;
    // rom_array[30814] = 32'hFFFFFFF1;
    // rom_array[30815] = 32'hFFFFFFF1;
    // rom_array[30816] = 32'hFFFFFFF1;
    // rom_array[30817] = 32'hFFFFFFF1;
    // rom_array[30818] = 32'hFFFFFFF1;
    // rom_array[30819] = 32'hFFFFFFF1;
    // rom_array[30820] = 32'hFFFFFFF1;
    // rom_array[30821] = 32'hFFFFFFF1;
    // rom_array[30822] = 32'hFFFFFFF1;
    // rom_array[30823] = 32'hFFFFFFF1;
    // rom_array[30824] = 32'hFFFFFFF1;
    // rom_array[30825] = 32'hFFFFFFF0;
    // rom_array[30826] = 32'hFFFFFFF0;
    // rom_array[30827] = 32'hFFFFFFF1;
    // rom_array[30828] = 32'hFFFFFFF1;
    // rom_array[30829] = 32'hFFFFFFF0;
    // rom_array[30830] = 32'hFFFFFFF0;
    // rom_array[30831] = 32'hFFFFFFF1;
    // rom_array[30832] = 32'hFFFFFFF1;
    // rom_array[30833] = 32'hFFFFFFF0;
    // rom_array[30834] = 32'hFFFFFFF0;
    // rom_array[30835] = 32'hFFFFFFF1;
    // rom_array[30836] = 32'hFFFFFFF1;
    // rom_array[30837] = 32'hFFFFFFF0;
    // rom_array[30838] = 32'hFFFFFFF0;
    // rom_array[30839] = 32'hFFFFFFF1;
    // rom_array[30840] = 32'hFFFFFFF1;
    // rom_array[30841] = 32'hFFFFFFF1;
    // rom_array[30842] = 32'hFFFFFFF1;
    // rom_array[30843] = 32'hFFFFFFF1;
    // rom_array[30844] = 32'hFFFFFFF1;
    // rom_array[30845] = 32'hFFFFFFF1;
    // rom_array[30846] = 32'hFFFFFFF1;
    // rom_array[30847] = 32'hFFFFFFF1;
    // rom_array[30848] = 32'hFFFFFFF1;
    // rom_array[30849] = 32'hFFFFFFF1;
    // rom_array[30850] = 32'hFFFFFFF1;
    // rom_array[30851] = 32'hFFFFFFF1;
    // rom_array[30852] = 32'hFFFFFFF1;
    // rom_array[30853] = 32'hFFFFFFF1;
    // rom_array[30854] = 32'hFFFFFFF1;
    // rom_array[30855] = 32'hFFFFFFF1;
    // rom_array[30856] = 32'hFFFFFFF1;
    // rom_array[30857] = 32'hFFFFFFF1;
    // rom_array[30858] = 32'hFFFFFFF1;
    // rom_array[30859] = 32'hFFFFFFF0;
    // rom_array[30860] = 32'hFFFFFFF0;
    // rom_array[30861] = 32'hFFFFFFF1;
    // rom_array[30862] = 32'hFFFFFFF1;
    // rom_array[30863] = 32'hFFFFFFF0;
    // rom_array[30864] = 32'hFFFFFFF0;
    // rom_array[30865] = 32'hFFFFFFF1;
    // rom_array[30866] = 32'hFFFFFFF1;
    // rom_array[30867] = 32'hFFFFFFF0;
    // rom_array[30868] = 32'hFFFFFFF0;
    // rom_array[30869] = 32'hFFFFFFF1;
    // rom_array[30870] = 32'hFFFFFFF1;
    // rom_array[30871] = 32'hFFFFFFF0;
    // rom_array[30872] = 32'hFFFFFFF0;
    // rom_array[30873] = 32'hFFFFFFF1;
    // rom_array[30874] = 32'hFFFFFFF1;
    // rom_array[30875] = 32'hFFFFFFF0;
    // rom_array[30876] = 32'hFFFFFFF0;
    // rom_array[30877] = 32'hFFFFFFF1;
    // rom_array[30878] = 32'hFFFFFFF1;
    // rom_array[30879] = 32'hFFFFFFF0;
    // rom_array[30880] = 32'hFFFFFFF0;
    // rom_array[30881] = 32'hFFFFFFF1;
    // rom_array[30882] = 32'hFFFFFFF1;
    // rom_array[30883] = 32'hFFFFFFF0;
    // rom_array[30884] = 32'hFFFFFFF0;
    // rom_array[30885] = 32'hFFFFFFF1;
    // rom_array[30886] = 32'hFFFFFFF1;
    // rom_array[30887] = 32'hFFFFFFF0;
    // rom_array[30888] = 32'hFFFFFFF0;
    // rom_array[30889] = 32'hFFFFFFF0;
    // rom_array[30890] = 32'hFFFFFFF0;
    // rom_array[30891] = 32'hFFFFFFF1;
    // rom_array[30892] = 32'hFFFFFFF1;
    // rom_array[30893] = 32'hFFFFFFF0;
    // rom_array[30894] = 32'hFFFFFFF0;
    // rom_array[30895] = 32'hFFFFFFF1;
    // rom_array[30896] = 32'hFFFFFFF1;
    // rom_array[30897] = 32'hFFFFFFF0;
    // rom_array[30898] = 32'hFFFFFFF0;
    // rom_array[30899] = 32'hFFFFFFF1;
    // rom_array[30900] = 32'hFFFFFFF1;
    // rom_array[30901] = 32'hFFFFFFF0;
    // rom_array[30902] = 32'hFFFFFFF0;
    // rom_array[30903] = 32'hFFFFFFF1;
    // rom_array[30904] = 32'hFFFFFFF1;
    // rom_array[30905] = 32'hFFFFFFF0;
    // rom_array[30906] = 32'hFFFFFFF0;
    // rom_array[30907] = 32'hFFFFFFF1;
    // rom_array[30908] = 32'hFFFFFFF1;
    // rom_array[30909] = 32'hFFFFFFF0;
    // rom_array[30910] = 32'hFFFFFFF0;
    // rom_array[30911] = 32'hFFFFFFF1;
    // rom_array[30912] = 32'hFFFFFFF1;
    // rom_array[30913] = 32'hFFFFFFF0;
    // rom_array[30914] = 32'hFFFFFFF0;
    // rom_array[30915] = 32'hFFFFFFF1;
    // rom_array[30916] = 32'hFFFFFFF1;
    // rom_array[30917] = 32'hFFFFFFF0;
    // rom_array[30918] = 32'hFFFFFFF0;
    // rom_array[30919] = 32'hFFFFFFF1;
    // rom_array[30920] = 32'hFFFFFFF1;
    // rom_array[30921] = 32'hFFFFFFF1;
    // rom_array[30922] = 32'hFFFFFFF1;
    // rom_array[30923] = 32'hFFFFFFF0;
    // rom_array[30924] = 32'hFFFFFFF0;
    // rom_array[30925] = 32'hFFFFFFF1;
    // rom_array[30926] = 32'hFFFFFFF1;
    // rom_array[30927] = 32'hFFFFFFF0;
    // rom_array[30928] = 32'hFFFFFFF0;
    // rom_array[30929] = 32'hFFFFFFF1;
    // rom_array[30930] = 32'hFFFFFFF1;
    // rom_array[30931] = 32'hFFFFFFF0;
    // rom_array[30932] = 32'hFFFFFFF0;
    // rom_array[30933] = 32'hFFFFFFF1;
    // rom_array[30934] = 32'hFFFFFFF1;
    // rom_array[30935] = 32'hFFFFFFF0;
    // rom_array[30936] = 32'hFFFFFFF0;
    // rom_array[30937] = 32'hFFFFFFF1;
    // rom_array[30938] = 32'hFFFFFFF1;
    // rom_array[30939] = 32'hFFFFFFF0;
    // rom_array[30940] = 32'hFFFFFFF0;
    // rom_array[30941] = 32'hFFFFFFF1;
    // rom_array[30942] = 32'hFFFFFFF1;
    // rom_array[30943] = 32'hFFFFFFF1;
    // rom_array[30944] = 32'hFFFFFFF1;
    // rom_array[30945] = 32'hFFFFFFF1;
    // rom_array[30946] = 32'hFFFFFFF1;
    // rom_array[30947] = 32'hFFFFFFF0;
    // rom_array[30948] = 32'hFFFFFFF0;
    // rom_array[30949] = 32'hFFFFFFF1;
    // rom_array[30950] = 32'hFFFFFFF1;
    // rom_array[30951] = 32'hFFFFFFF1;
    // rom_array[30952] = 32'hFFFFFFF1;
    // rom_array[30953] = 32'hFFFFFFF0;
    // rom_array[30954] = 32'hFFFFFFF0;
    // rom_array[30955] = 32'hFFFFFFF1;
    // rom_array[30956] = 32'hFFFFFFF1;
    // rom_array[30957] = 32'hFFFFFFF0;
    // rom_array[30958] = 32'hFFFFFFF0;
    // rom_array[30959] = 32'hFFFFFFF0;
    // rom_array[30960] = 32'hFFFFFFF0;
    // rom_array[30961] = 32'hFFFFFFF0;
    // rom_array[30962] = 32'hFFFFFFF0;
    // rom_array[30963] = 32'hFFFFFFF1;
    // rom_array[30964] = 32'hFFFFFFF1;
    // rom_array[30965] = 32'hFFFFFFF0;
    // rom_array[30966] = 32'hFFFFFFF0;
    // rom_array[30967] = 32'hFFFFFFF0;
    // rom_array[30968] = 32'hFFFFFFF0;
    // rom_array[30969] = 32'hFFFFFFF1;
    // rom_array[30970] = 32'hFFFFFFF1;
    // rom_array[30971] = 32'hFFFFFFF1;
    // rom_array[30972] = 32'hFFFFFFF1;
    // rom_array[30973] = 32'hFFFFFFF0;
    // rom_array[30974] = 32'hFFFFFFF0;
    // rom_array[30975] = 32'hFFFFFFF0;
    // rom_array[30976] = 32'hFFFFFFF0;
    // rom_array[30977] = 32'hFFFFFFF1;
    // rom_array[30978] = 32'hFFFFFFF1;
    // rom_array[30979] = 32'hFFFFFFF1;
    // rom_array[30980] = 32'hFFFFFFF1;
    // rom_array[30981] = 32'hFFFFFFF0;
    // rom_array[30982] = 32'hFFFFFFF0;
    // rom_array[30983] = 32'hFFFFFFF0;
    // rom_array[30984] = 32'hFFFFFFF0;
    // rom_array[30985] = 32'hFFFFFFF1;
    // rom_array[30986] = 32'hFFFFFFF1;
    // rom_array[30987] = 32'hFFFFFFF1;
    // rom_array[30988] = 32'hFFFFFFF1;
    // rom_array[30989] = 32'hFFFFFFF0;
    // rom_array[30990] = 32'hFFFFFFF0;
    // rom_array[30991] = 32'hFFFFFFF0;
    // rom_array[30992] = 32'hFFFFFFF0;
    // rom_array[30993] = 32'hFFFFFFF1;
    // rom_array[30994] = 32'hFFFFFFF1;
    // rom_array[30995] = 32'hFFFFFFF1;
    // rom_array[30996] = 32'hFFFFFFF1;
    // rom_array[30997] = 32'hFFFFFFF0;
    // rom_array[30998] = 32'hFFFFFFF0;
    // rom_array[30999] = 32'hFFFFFFF0;
    // rom_array[31000] = 32'hFFFFFFF0;
    // rom_array[31001] = 32'hFFFFFFF1;
    // rom_array[31002] = 32'hFFFFFFF1;
    // rom_array[31003] = 32'hFFFFFFF1;
    // rom_array[31004] = 32'hFFFFFFF1;
    // rom_array[31005] = 32'hFFFFFFF1;
    // rom_array[31006] = 32'hFFFFFFF1;
    // rom_array[31007] = 32'hFFFFFFF1;
    // rom_array[31008] = 32'hFFFFFFF1;
    // rom_array[31009] = 32'hFFFFFFF1;
    // rom_array[31010] = 32'hFFFFFFF1;
    // rom_array[31011] = 32'hFFFFFFF1;
    // rom_array[31012] = 32'hFFFFFFF1;
    // rom_array[31013] = 32'hFFFFFFF1;
    // rom_array[31014] = 32'hFFFFFFF1;
    // rom_array[31015] = 32'hFFFFFFF1;
    // rom_array[31016] = 32'hFFFFFFF1;
    // rom_array[31017] = 32'hFFFFFFF1;
    // rom_array[31018] = 32'hFFFFFFF1;
    // rom_array[31019] = 32'hFFFFFFF1;
    // rom_array[31020] = 32'hFFFFFFF1;
    // rom_array[31021] = 32'hFFFFFFF1;
    // rom_array[31022] = 32'hFFFFFFF1;
    // rom_array[31023] = 32'hFFFFFFF1;
    // rom_array[31024] = 32'hFFFFFFF1;
    // rom_array[31025] = 32'hFFFFFFF1;
    // rom_array[31026] = 32'hFFFFFFF1;
    // rom_array[31027] = 32'hFFFFFFF1;
    // rom_array[31028] = 32'hFFFFFFF1;
    // rom_array[31029] = 32'hFFFFFFF1;
    // rom_array[31030] = 32'hFFFFFFF1;
    // rom_array[31031] = 32'hFFFFFFF1;
    // rom_array[31032] = 32'hFFFFFFF1;
    // rom_array[31033] = 32'hFFFFFFF0;
    // rom_array[31034] = 32'hFFFFFFF0;
    // rom_array[31035] = 32'hFFFFFFF1;
    // rom_array[31036] = 32'hFFFFFFF1;
    // rom_array[31037] = 32'hFFFFFFF0;
    // rom_array[31038] = 32'hFFFFFFF0;
    // rom_array[31039] = 32'hFFFFFFF1;
    // rom_array[31040] = 32'hFFFFFFF1;
    // rom_array[31041] = 32'hFFFFFFF0;
    // rom_array[31042] = 32'hFFFFFFF0;
    // rom_array[31043] = 32'hFFFFFFF1;
    // rom_array[31044] = 32'hFFFFFFF1;
    // rom_array[31045] = 32'hFFFFFFF0;
    // rom_array[31046] = 32'hFFFFFFF0;
    // rom_array[31047] = 32'hFFFFFFF1;
    // rom_array[31048] = 32'hFFFFFFF1;
    // rom_array[31049] = 32'hFFFFFFF1;
    // rom_array[31050] = 32'hFFFFFFF1;
    // rom_array[31051] = 32'hFFFFFFF1;
    // rom_array[31052] = 32'hFFFFFFF1;
    // rom_array[31053] = 32'hFFFFFFF1;
    // rom_array[31054] = 32'hFFFFFFF1;
    // rom_array[31055] = 32'hFFFFFFF1;
    // rom_array[31056] = 32'hFFFFFFF1;
    // rom_array[31057] = 32'hFFFFFFF1;
    // rom_array[31058] = 32'hFFFFFFF1;
    // rom_array[31059] = 32'hFFFFFFF1;
    // rom_array[31060] = 32'hFFFFFFF1;
    // rom_array[31061] = 32'hFFFFFFF1;
    // rom_array[31062] = 32'hFFFFFFF1;
    // rom_array[31063] = 32'hFFFFFFF1;
    // rom_array[31064] = 32'hFFFFFFF1;
    // rom_array[31065] = 32'hFFFFFFF0;
    // rom_array[31066] = 32'hFFFFFFF0;
    // rom_array[31067] = 32'hFFFFFFF1;
    // rom_array[31068] = 32'hFFFFFFF1;
    // rom_array[31069] = 32'hFFFFFFF0;
    // rom_array[31070] = 32'hFFFFFFF0;
    // rom_array[31071] = 32'hFFFFFFF0;
    // rom_array[31072] = 32'hFFFFFFF0;
    // rom_array[31073] = 32'hFFFFFFF0;
    // rom_array[31074] = 32'hFFFFFFF0;
    // rom_array[31075] = 32'hFFFFFFF1;
    // rom_array[31076] = 32'hFFFFFFF1;
    // rom_array[31077] = 32'hFFFFFFF0;
    // rom_array[31078] = 32'hFFFFFFF0;
    // rom_array[31079] = 32'hFFFFFFF0;
    // rom_array[31080] = 32'hFFFFFFF0;
    // rom_array[31081] = 32'hFFFFFFF1;
    // rom_array[31082] = 32'hFFFFFFF1;
    // rom_array[31083] = 32'hFFFFFFF1;
    // rom_array[31084] = 32'hFFFFFFF1;
    // rom_array[31085] = 32'hFFFFFFF0;
    // rom_array[31086] = 32'hFFFFFFF0;
    // rom_array[31087] = 32'hFFFFFFF0;
    // rom_array[31088] = 32'hFFFFFFF0;
    // rom_array[31089] = 32'hFFFFFFF1;
    // rom_array[31090] = 32'hFFFFFFF1;
    // rom_array[31091] = 32'hFFFFFFF1;
    // rom_array[31092] = 32'hFFFFFFF1;
    // rom_array[31093] = 32'hFFFFFFF0;
    // rom_array[31094] = 32'hFFFFFFF0;
    // rom_array[31095] = 32'hFFFFFFF0;
    // rom_array[31096] = 32'hFFFFFFF0;
    // rom_array[31097] = 32'hFFFFFFF1;
    // rom_array[31098] = 32'hFFFFFFF1;
    // rom_array[31099] = 32'hFFFFFFF1;
    // rom_array[31100] = 32'hFFFFFFF1;
    // rom_array[31101] = 32'hFFFFFFF1;
    // rom_array[31102] = 32'hFFFFFFF1;
    // rom_array[31103] = 32'hFFFFFFF1;
    // rom_array[31104] = 32'hFFFFFFF1;
    // rom_array[31105] = 32'hFFFFFFF1;
    // rom_array[31106] = 32'hFFFFFFF1;
    // rom_array[31107] = 32'hFFFFFFF1;
    // rom_array[31108] = 32'hFFFFFFF1;
    // rom_array[31109] = 32'hFFFFFFF1;
    // rom_array[31110] = 32'hFFFFFFF1;
    // rom_array[31111] = 32'hFFFFFFF1;
    // rom_array[31112] = 32'hFFFFFFF1;
    // rom_array[31113] = 32'hFFFFFFF1;
    // rom_array[31114] = 32'hFFFFFFF1;
    // rom_array[31115] = 32'hFFFFFFF1;
    // rom_array[31116] = 32'hFFFFFFF1;
    // rom_array[31117] = 32'hFFFFFFF0;
    // rom_array[31118] = 32'hFFFFFFF0;
    // rom_array[31119] = 32'hFFFFFFF0;
    // rom_array[31120] = 32'hFFFFFFF0;
    // rom_array[31121] = 32'hFFFFFFF1;
    // rom_array[31122] = 32'hFFFFFFF1;
    // rom_array[31123] = 32'hFFFFFFF1;
    // rom_array[31124] = 32'hFFFFFFF1;
    // rom_array[31125] = 32'hFFFFFFF0;
    // rom_array[31126] = 32'hFFFFFFF0;
    // rom_array[31127] = 32'hFFFFFFF0;
    // rom_array[31128] = 32'hFFFFFFF0;
    // rom_array[31129] = 32'hFFFFFFF1;
    // rom_array[31130] = 32'hFFFFFFF1;
    // rom_array[31131] = 32'hFFFFFFF1;
    // rom_array[31132] = 32'hFFFFFFF1;
    // rom_array[31133] = 32'hFFFFFFF0;
    // rom_array[31134] = 32'hFFFFFFF0;
    // rom_array[31135] = 32'hFFFFFFF0;
    // rom_array[31136] = 32'hFFFFFFF0;
    // rom_array[31137] = 32'hFFFFFFF1;
    // rom_array[31138] = 32'hFFFFFFF1;
    // rom_array[31139] = 32'hFFFFFFF1;
    // rom_array[31140] = 32'hFFFFFFF1;
    // rom_array[31141] = 32'hFFFFFFF0;
    // rom_array[31142] = 32'hFFFFFFF0;
    // rom_array[31143] = 32'hFFFFFFF0;
    // rom_array[31144] = 32'hFFFFFFF0;
    // rom_array[31145] = 32'hFFFFFFF1;
    // rom_array[31146] = 32'hFFFFFFF1;
    // rom_array[31147] = 32'hFFFFFFF1;
    // rom_array[31148] = 32'hFFFFFFF1;
    // rom_array[31149] = 32'hFFFFFFF0;
    // rom_array[31150] = 32'hFFFFFFF0;
    // rom_array[31151] = 32'hFFFFFFF0;
    // rom_array[31152] = 32'hFFFFFFF0;
    // rom_array[31153] = 32'hFFFFFFF1;
    // rom_array[31154] = 32'hFFFFFFF1;
    // rom_array[31155] = 32'hFFFFFFF1;
    // rom_array[31156] = 32'hFFFFFFF1;
    // rom_array[31157] = 32'hFFFFFFF0;
    // rom_array[31158] = 32'hFFFFFFF0;
    // rom_array[31159] = 32'hFFFFFFF0;
    // rom_array[31160] = 32'hFFFFFFF0;
    // rom_array[31161] = 32'hFFFFFFF1;
    // rom_array[31162] = 32'hFFFFFFF1;
    // rom_array[31163] = 32'hFFFFFFF1;
    // rom_array[31164] = 32'hFFFFFFF1;
    // rom_array[31165] = 32'hFFFFFFF0;
    // rom_array[31166] = 32'hFFFFFFF0;
    // rom_array[31167] = 32'hFFFFFFF0;
    // rom_array[31168] = 32'hFFFFFFF0;
    // rom_array[31169] = 32'hFFFFFFF1;
    // rom_array[31170] = 32'hFFFFFFF1;
    // rom_array[31171] = 32'hFFFFFFF1;
    // rom_array[31172] = 32'hFFFFFFF1;
    // rom_array[31173] = 32'hFFFFFFF0;
    // rom_array[31174] = 32'hFFFFFFF0;
    // rom_array[31175] = 32'hFFFFFFF0;
    // rom_array[31176] = 32'hFFFFFFF0;
    // rom_array[31177] = 32'hFFFFFFF1;
    // rom_array[31178] = 32'hFFFFFFF1;
    // rom_array[31179] = 32'hFFFFFFF1;
    // rom_array[31180] = 32'hFFFFFFF1;
    // rom_array[31181] = 32'hFFFFFFF0;
    // rom_array[31182] = 32'hFFFFFFF0;
    // rom_array[31183] = 32'hFFFFFFF0;
    // rom_array[31184] = 32'hFFFFFFF0;
    // rom_array[31185] = 32'hFFFFFFF1;
    // rom_array[31186] = 32'hFFFFFFF1;
    // rom_array[31187] = 32'hFFFFFFF1;
    // rom_array[31188] = 32'hFFFFFFF1;
    // rom_array[31189] = 32'hFFFFFFF0;
    // rom_array[31190] = 32'hFFFFFFF0;
    // rom_array[31191] = 32'hFFFFFFF0;
    // rom_array[31192] = 32'hFFFFFFF0;
    // rom_array[31193] = 32'hFFFFFFF1;
    // rom_array[31194] = 32'hFFFFFFF1;
    // rom_array[31195] = 32'hFFFFFFF1;
    // rom_array[31196] = 32'hFFFFFFF1;
    // rom_array[31197] = 32'hFFFFFFF0;
    // rom_array[31198] = 32'hFFFFFFF0;
    // rom_array[31199] = 32'hFFFFFFF0;
    // rom_array[31200] = 32'hFFFFFFF0;
    // rom_array[31201] = 32'hFFFFFFF1;
    // rom_array[31202] = 32'hFFFFFFF1;
    // rom_array[31203] = 32'hFFFFFFF1;
    // rom_array[31204] = 32'hFFFFFFF1;
    // rom_array[31205] = 32'hFFFFFFF0;
    // rom_array[31206] = 32'hFFFFFFF0;
    // rom_array[31207] = 32'hFFFFFFF0;
    // rom_array[31208] = 32'hFFFFFFF0;
    // rom_array[31209] = 32'hFFFFFFF1;
    // rom_array[31210] = 32'hFFFFFFF1;
    // rom_array[31211] = 32'hFFFFFFF1;
    // rom_array[31212] = 32'hFFFFFFF1;
    // rom_array[31213] = 32'hFFFFFFF0;
    // rom_array[31214] = 32'hFFFFFFF0;
    // rom_array[31215] = 32'hFFFFFFF0;
    // rom_array[31216] = 32'hFFFFFFF0;
    // rom_array[31217] = 32'hFFFFFFF1;
    // rom_array[31218] = 32'hFFFFFFF1;
    // rom_array[31219] = 32'hFFFFFFF1;
    // rom_array[31220] = 32'hFFFFFFF1;
    // rom_array[31221] = 32'hFFFFFFF0;
    // rom_array[31222] = 32'hFFFFFFF0;
    // rom_array[31223] = 32'hFFFFFFF0;
    // rom_array[31224] = 32'hFFFFFFF0;
    // rom_array[31225] = 32'hFFFFFFF1;
    // rom_array[31226] = 32'hFFFFFFF1;
    // rom_array[31227] = 32'hFFFFFFF1;
    // rom_array[31228] = 32'hFFFFFFF1;
    // rom_array[31229] = 32'hFFFFFFF0;
    // rom_array[31230] = 32'hFFFFFFF0;
    // rom_array[31231] = 32'hFFFFFFF0;
    // rom_array[31232] = 32'hFFFFFFF0;
    // rom_array[31233] = 32'hFFFFFFF1;
    // rom_array[31234] = 32'hFFFFFFF1;
    // rom_array[31235] = 32'hFFFFFFF1;
    // rom_array[31236] = 32'hFFFFFFF1;
    // rom_array[31237] = 32'hFFFFFFF0;
    // rom_array[31238] = 32'hFFFFFFF0;
    // rom_array[31239] = 32'hFFFFFFF0;
    // rom_array[31240] = 32'hFFFFFFF0;
    // rom_array[31241] = 32'hFFFFFFF1;
    // rom_array[31242] = 32'hFFFFFFF1;
    // rom_array[31243] = 32'hFFFFFFF1;
    // rom_array[31244] = 32'hFFFFFFF1;
    // rom_array[31245] = 32'hFFFFFFF1;
    // rom_array[31246] = 32'hFFFFFFF1;
    // rom_array[31247] = 32'hFFFFFFF1;
    // rom_array[31248] = 32'hFFFFFFF1;
    // rom_array[31249] = 32'hFFFFFFF1;
    // rom_array[31250] = 32'hFFFFFFF1;
    // rom_array[31251] = 32'hFFFFFFF1;
    // rom_array[31252] = 32'hFFFFFFF1;
    // rom_array[31253] = 32'hFFFFFFF1;
    // rom_array[31254] = 32'hFFFFFFF1;
    // rom_array[31255] = 32'hFFFFFFF1;
    // rom_array[31256] = 32'hFFFFFFF1;
    // rom_array[31257] = 32'hFFFFFFF1;
    // rom_array[31258] = 32'hFFFFFFF1;
    // rom_array[31259] = 32'hFFFFFFF1;
    // rom_array[31260] = 32'hFFFFFFF1;
    // rom_array[31261] = 32'hFFFFFFF0;
    // rom_array[31262] = 32'hFFFFFFF0;
    // rom_array[31263] = 32'hFFFFFFF0;
    // rom_array[31264] = 32'hFFFFFFF0;
    // rom_array[31265] = 32'hFFFFFFF1;
    // rom_array[31266] = 32'hFFFFFFF1;
    // rom_array[31267] = 32'hFFFFFFF1;
    // rom_array[31268] = 32'hFFFFFFF1;
    // rom_array[31269] = 32'hFFFFFFF0;
    // rom_array[31270] = 32'hFFFFFFF0;
    // rom_array[31271] = 32'hFFFFFFF0;
    // rom_array[31272] = 32'hFFFFFFF0;
    // rom_array[31273] = 32'hFFFFFFF1;
    // rom_array[31274] = 32'hFFFFFFF1;
    // rom_array[31275] = 32'hFFFFFFF1;
    // rom_array[31276] = 32'hFFFFFFF1;
    // rom_array[31277] = 32'hFFFFFFF0;
    // rom_array[31278] = 32'hFFFFFFF0;
    // rom_array[31279] = 32'hFFFFFFF0;
    // rom_array[31280] = 32'hFFFFFFF0;
    // rom_array[31281] = 32'hFFFFFFF1;
    // rom_array[31282] = 32'hFFFFFFF1;
    // rom_array[31283] = 32'hFFFFFFF1;
    // rom_array[31284] = 32'hFFFFFFF1;
    // rom_array[31285] = 32'hFFFFFFF0;
    // rom_array[31286] = 32'hFFFFFFF0;
    // rom_array[31287] = 32'hFFFFFFF0;
    // rom_array[31288] = 32'hFFFFFFF0;
    // rom_array[31289] = 32'hFFFFFFF0;
    // rom_array[31290] = 32'hFFFFFFF0;
    // rom_array[31291] = 32'hFFFFFFF0;
    // rom_array[31292] = 32'hFFFFFFF0;
    // rom_array[31293] = 32'hFFFFFFF0;
    // rom_array[31294] = 32'hFFFFFFF0;
    // rom_array[31295] = 32'hFFFFFFF1;
    // rom_array[31296] = 32'hFFFFFFF1;
    // rom_array[31297] = 32'hFFFFFFF0;
    // rom_array[31298] = 32'hFFFFFFF0;
    // rom_array[31299] = 32'hFFFFFFF0;
    // rom_array[31300] = 32'hFFFFFFF0;
    // rom_array[31301] = 32'hFFFFFFF0;
    // rom_array[31302] = 32'hFFFFFFF0;
    // rom_array[31303] = 32'hFFFFFFF1;
    // rom_array[31304] = 32'hFFFFFFF1;
    // rom_array[31305] = 32'hFFFFFFF0;
    // rom_array[31306] = 32'hFFFFFFF0;
    // rom_array[31307] = 32'hFFFFFFF0;
    // rom_array[31308] = 32'hFFFFFFF0;
    // rom_array[31309] = 32'hFFFFFFF1;
    // rom_array[31310] = 32'hFFFFFFF1;
    // rom_array[31311] = 32'hFFFFFFF1;
    // rom_array[31312] = 32'hFFFFFFF1;
    // rom_array[31313] = 32'hFFFFFFF0;
    // rom_array[31314] = 32'hFFFFFFF0;
    // rom_array[31315] = 32'hFFFFFFF0;
    // rom_array[31316] = 32'hFFFFFFF0;
    // rom_array[31317] = 32'hFFFFFFF1;
    // rom_array[31318] = 32'hFFFFFFF1;
    // rom_array[31319] = 32'hFFFFFFF1;
    // rom_array[31320] = 32'hFFFFFFF1;
    // rom_array[31321] = 32'hFFFFFFF0;
    // rom_array[31322] = 32'hFFFFFFF0;
    // rom_array[31323] = 32'hFFFFFFF0;
    // rom_array[31324] = 32'hFFFFFFF0;
    // rom_array[31325] = 32'hFFFFFFF1;
    // rom_array[31326] = 32'hFFFFFFF1;
    // rom_array[31327] = 32'hFFFFFFF1;
    // rom_array[31328] = 32'hFFFFFFF1;
    // rom_array[31329] = 32'hFFFFFFF0;
    // rom_array[31330] = 32'hFFFFFFF0;
    // rom_array[31331] = 32'hFFFFFFF0;
    // rom_array[31332] = 32'hFFFFFFF0;
    // rom_array[31333] = 32'hFFFFFFF1;
    // rom_array[31334] = 32'hFFFFFFF1;
    // rom_array[31335] = 32'hFFFFFFF1;
    // rom_array[31336] = 32'hFFFFFFF1;
    // rom_array[31337] = 32'hFFFFFFF0;
    // rom_array[31338] = 32'hFFFFFFF0;
    // rom_array[31339] = 32'hFFFFFFF0;
    // rom_array[31340] = 32'hFFFFFFF0;
    // rom_array[31341] = 32'hFFFFFFF1;
    // rom_array[31342] = 32'hFFFFFFF1;
    // rom_array[31343] = 32'hFFFFFFF1;
    // rom_array[31344] = 32'hFFFFFFF1;
    // rom_array[31345] = 32'hFFFFFFF0;
    // rom_array[31346] = 32'hFFFFFFF0;
    // rom_array[31347] = 32'hFFFFFFF0;
    // rom_array[31348] = 32'hFFFFFFF0;
    // rom_array[31349] = 32'hFFFFFFF1;
    // rom_array[31350] = 32'hFFFFFFF1;
    // rom_array[31351] = 32'hFFFFFFF1;
    // rom_array[31352] = 32'hFFFFFFF1;
    // rom_array[31353] = 32'hFFFFFFF0;
    // rom_array[31354] = 32'hFFFFFFF0;
    // rom_array[31355] = 32'hFFFFFFF1;
    // rom_array[31356] = 32'hFFFFFFF1;
    // rom_array[31357] = 32'hFFFFFFF0;
    // rom_array[31358] = 32'hFFFFFFF0;
    // rom_array[31359] = 32'hFFFFFFF1;
    // rom_array[31360] = 32'hFFFFFFF1;
    // rom_array[31361] = 32'hFFFFFFF0;
    // rom_array[31362] = 32'hFFFFFFF0;
    // rom_array[31363] = 32'hFFFFFFF1;
    // rom_array[31364] = 32'hFFFFFFF1;
    // rom_array[31365] = 32'hFFFFFFF0;
    // rom_array[31366] = 32'hFFFFFFF0;
    // rom_array[31367] = 32'hFFFFFFF1;
    // rom_array[31368] = 32'hFFFFFFF1;
    // rom_array[31369] = 32'hFFFFFFF0;
    // rom_array[31370] = 32'hFFFFFFF0;
    // rom_array[31371] = 32'hFFFFFFF1;
    // rom_array[31372] = 32'hFFFFFFF1;
    // rom_array[31373] = 32'hFFFFFFF0;
    // rom_array[31374] = 32'hFFFFFFF0;
    // rom_array[31375] = 32'hFFFFFFF1;
    // rom_array[31376] = 32'hFFFFFFF1;
    // rom_array[31377] = 32'hFFFFFFF0;
    // rom_array[31378] = 32'hFFFFFFF0;
    // rom_array[31379] = 32'hFFFFFFF1;
    // rom_array[31380] = 32'hFFFFFFF1;
    // rom_array[31381] = 32'hFFFFFFF0;
    // rom_array[31382] = 32'hFFFFFFF0;
    // rom_array[31383] = 32'hFFFFFFF1;
    // rom_array[31384] = 32'hFFFFFFF1;
    // rom_array[31385] = 32'hFFFFFFF0;
    // rom_array[31386] = 32'hFFFFFFF0;
    // rom_array[31387] = 32'hFFFFFFF1;
    // rom_array[31388] = 32'hFFFFFFF1;
    // rom_array[31389] = 32'hFFFFFFF0;
    // rom_array[31390] = 32'hFFFFFFF0;
    // rom_array[31391] = 32'hFFFFFFF1;
    // rom_array[31392] = 32'hFFFFFFF1;
    // rom_array[31393] = 32'hFFFFFFF0;
    // rom_array[31394] = 32'hFFFFFFF0;
    // rom_array[31395] = 32'hFFFFFFF1;
    // rom_array[31396] = 32'hFFFFFFF1;
    // rom_array[31397] = 32'hFFFFFFF0;
    // rom_array[31398] = 32'hFFFFFFF0;
    // rom_array[31399] = 32'hFFFFFFF1;
    // rom_array[31400] = 32'hFFFFFFF1;
    // rom_array[31401] = 32'hFFFFFFF0;
    // rom_array[31402] = 32'hFFFFFFF0;
    // rom_array[31403] = 32'hFFFFFFF1;
    // rom_array[31404] = 32'hFFFFFFF1;
    // rom_array[31405] = 32'hFFFFFFF0;
    // rom_array[31406] = 32'hFFFFFFF0;
    // rom_array[31407] = 32'hFFFFFFF1;
    // rom_array[31408] = 32'hFFFFFFF1;
    // rom_array[31409] = 32'hFFFFFFF0;
    // rom_array[31410] = 32'hFFFFFFF0;
    // rom_array[31411] = 32'hFFFFFFF1;
    // rom_array[31412] = 32'hFFFFFFF1;
    // rom_array[31413] = 32'hFFFFFFF0;
    // rom_array[31414] = 32'hFFFFFFF0;
    // rom_array[31415] = 32'hFFFFFFF1;
    // rom_array[31416] = 32'hFFFFFFF1;
    // rom_array[31417] = 32'hFFFFFFF0;
    // rom_array[31418] = 32'hFFFFFFF0;
    // rom_array[31419] = 32'hFFFFFFF1;
    // rom_array[31420] = 32'hFFFFFFF1;
    // rom_array[31421] = 32'hFFFFFFF0;
    // rom_array[31422] = 32'hFFFFFFF0;
    // rom_array[31423] = 32'hFFFFFFF1;
    // rom_array[31424] = 32'hFFFFFFF1;
    // rom_array[31425] = 32'hFFFFFFF0;
    // rom_array[31426] = 32'hFFFFFFF0;
    // rom_array[31427] = 32'hFFFFFFF1;
    // rom_array[31428] = 32'hFFFFFFF1;
    // rom_array[31429] = 32'hFFFFFFF0;
    // rom_array[31430] = 32'hFFFFFFF0;
    // rom_array[31431] = 32'hFFFFFFF1;
    // rom_array[31432] = 32'hFFFFFFF1;
    // rom_array[31433] = 32'hFFFFFFF0;
    // rom_array[31434] = 32'hFFFFFFF0;
    // rom_array[31435] = 32'hFFFFFFF1;
    // rom_array[31436] = 32'hFFFFFFF1;
    // rom_array[31437] = 32'hFFFFFFF0;
    // rom_array[31438] = 32'hFFFFFFF0;
    // rom_array[31439] = 32'hFFFFFFF1;
    // rom_array[31440] = 32'hFFFFFFF1;
    // rom_array[31441] = 32'hFFFFFFF0;
    // rom_array[31442] = 32'hFFFFFFF0;
    // rom_array[31443] = 32'hFFFFFFF1;
    // rom_array[31444] = 32'hFFFFFFF1;
    // rom_array[31445] = 32'hFFFFFFF0;
    // rom_array[31446] = 32'hFFFFFFF0;
    // rom_array[31447] = 32'hFFFFFFF1;
    // rom_array[31448] = 32'hFFFFFFF1;
    // rom_array[31449] = 32'hFFFFFFF0;
    // rom_array[31450] = 32'hFFFFFFF0;
    // rom_array[31451] = 32'hFFFFFFF0;
    // rom_array[31452] = 32'hFFFFFFF0;
    // rom_array[31453] = 32'hFFFFFFF1;
    // rom_array[31454] = 32'hFFFFFFF1;
    // rom_array[31455] = 32'hFFFFFFF1;
    // rom_array[31456] = 32'hFFFFFFF1;
    // rom_array[31457] = 32'hFFFFFFF0;
    // rom_array[31458] = 32'hFFFFFFF0;
    // rom_array[31459] = 32'hFFFFFFF0;
    // rom_array[31460] = 32'hFFFFFFF0;
    // rom_array[31461] = 32'hFFFFFFF1;
    // rom_array[31462] = 32'hFFFFFFF1;
    // rom_array[31463] = 32'hFFFFFFF1;
    // rom_array[31464] = 32'hFFFFFFF1;
    // rom_array[31465] = 32'hFFFFFFF1;
    // rom_array[31466] = 32'hFFFFFFF1;
    // rom_array[31467] = 32'hFFFFFFF1;
    // rom_array[31468] = 32'hFFFFFFF1;
    // rom_array[31469] = 32'hFFFFFFF1;
    // rom_array[31470] = 32'hFFFFFFF1;
    // rom_array[31471] = 32'hFFFFFFF1;
    // rom_array[31472] = 32'hFFFFFFF1;
    // rom_array[31473] = 32'hFFFFFFF1;
    // rom_array[31474] = 32'hFFFFFFF1;
    // rom_array[31475] = 32'hFFFFFFF1;
    // rom_array[31476] = 32'hFFFFFFF1;
    // rom_array[31477] = 32'hFFFFFFF1;
    // rom_array[31478] = 32'hFFFFFFF1;
    // rom_array[31479] = 32'hFFFFFFF1;
    // rom_array[31480] = 32'hFFFFFFF1;
    // rom_array[31481] = 32'hFFFFFFF1;
    // rom_array[31482] = 32'hFFFFFFF1;
    // rom_array[31483] = 32'hFFFFFFF1;
    // rom_array[31484] = 32'hFFFFFFF1;
    // rom_array[31485] = 32'hFFFFFFF1;
    // rom_array[31486] = 32'hFFFFFFF1;
    // rom_array[31487] = 32'hFFFFFFF1;
    // rom_array[31488] = 32'hFFFFFFF1;
    // rom_array[31489] = 32'hFFFFFFF1;
    // rom_array[31490] = 32'hFFFFFFF1;
    // rom_array[31491] = 32'hFFFFFFF1;
    // rom_array[31492] = 32'hFFFFFFF1;
    // rom_array[31493] = 32'hFFFFFFF1;
    // rom_array[31494] = 32'hFFFFFFF1;
    // rom_array[31495] = 32'hFFFFFFF1;
    // rom_array[31496] = 32'hFFFFFFF1;
    // rom_array[31497] = 32'hFFFFFFF1;
    // rom_array[31498] = 32'hFFFFFFF1;
    // rom_array[31499] = 32'hFFFFFFF1;
    // rom_array[31500] = 32'hFFFFFFF1;
    // rom_array[31501] = 32'hFFFFFFF1;
    // rom_array[31502] = 32'hFFFFFFF1;
    // rom_array[31503] = 32'hFFFFFFF1;
    // rom_array[31504] = 32'hFFFFFFF1;
    // rom_array[31505] = 32'hFFFFFFF1;
    // rom_array[31506] = 32'hFFFFFFF1;
    // rom_array[31507] = 32'hFFFFFFF1;
    // rom_array[31508] = 32'hFFFFFFF1;
    // rom_array[31509] = 32'hFFFFFFF1;
    // rom_array[31510] = 32'hFFFFFFF1;
    // rom_array[31511] = 32'hFFFFFFF1;
    // rom_array[31512] = 32'hFFFFFFF1;
    // rom_array[31513] = 32'hFFFFFFF1;
    // rom_array[31514] = 32'hFFFFFFF1;
    // rom_array[31515] = 32'hFFFFFFF1;
    // rom_array[31516] = 32'hFFFFFFF1;
    // rom_array[31517] = 32'hFFFFFFF1;
    // rom_array[31518] = 32'hFFFFFFF1;
    // rom_array[31519] = 32'hFFFFFFF1;
    // rom_array[31520] = 32'hFFFFFFF1;
    // rom_array[31521] = 32'hFFFFFFF1;
    // rom_array[31522] = 32'hFFFFFFF1;
    // rom_array[31523] = 32'hFFFFFFF1;
    // rom_array[31524] = 32'hFFFFFFF1;
    // rom_array[31525] = 32'hFFFFFFF1;
    // rom_array[31526] = 32'hFFFFFFF1;
    // rom_array[31527] = 32'hFFFFFFF1;
    // rom_array[31528] = 32'hFFFFFFF1;
    // rom_array[31529] = 32'hFFFFFFF1;
    // rom_array[31530] = 32'hFFFFFFF1;
    // rom_array[31531] = 32'hFFFFFFF1;
    // rom_array[31532] = 32'hFFFFFFF1;
    // rom_array[31533] = 32'hFFFFFFF1;
    // rom_array[31534] = 32'hFFFFFFF1;
    // rom_array[31535] = 32'hFFFFFFF1;
    // rom_array[31536] = 32'hFFFFFFF1;
    // rom_array[31537] = 32'hFFFFFFF1;
    // rom_array[31538] = 32'hFFFFFFF1;
    // rom_array[31539] = 32'hFFFFFFF1;
    // rom_array[31540] = 32'hFFFFFFF1;
    // rom_array[31541] = 32'hFFFFFFF1;
    // rom_array[31542] = 32'hFFFFFFF1;
    // rom_array[31543] = 32'hFFFFFFF1;
    // rom_array[31544] = 32'hFFFFFFF1;
    // rom_array[31545] = 32'hFFFFFFF0;
    // rom_array[31546] = 32'hFFFFFFF0;
    // rom_array[31547] = 32'hFFFFFFF0;
    // rom_array[31548] = 32'hFFFFFFF0;
    // rom_array[31549] = 32'hFFFFFFF1;
    // rom_array[31550] = 32'hFFFFFFF1;
    // rom_array[31551] = 32'hFFFFFFF1;
    // rom_array[31552] = 32'hFFFFFFF1;
    // rom_array[31553] = 32'hFFFFFFF0;
    // rom_array[31554] = 32'hFFFFFFF0;
    // rom_array[31555] = 32'hFFFFFFF0;
    // rom_array[31556] = 32'hFFFFFFF0;
    // rom_array[31557] = 32'hFFFFFFF1;
    // rom_array[31558] = 32'hFFFFFFF1;
    // rom_array[31559] = 32'hFFFFFFF1;
    // rom_array[31560] = 32'hFFFFFFF1;
    // rom_array[31561] = 32'hFFFFFFF1;
    // rom_array[31562] = 32'hFFFFFFF1;
    // rom_array[31563] = 32'hFFFFFFF1;
    // rom_array[31564] = 32'hFFFFFFF1;
    // rom_array[31565] = 32'hFFFFFFF1;
    // rom_array[31566] = 32'hFFFFFFF1;
    // rom_array[31567] = 32'hFFFFFFF1;
    // rom_array[31568] = 32'hFFFFFFF1;
    // rom_array[31569] = 32'hFFFFFFF1;
    // rom_array[31570] = 32'hFFFFFFF1;
    // rom_array[31571] = 32'hFFFFFFF1;
    // rom_array[31572] = 32'hFFFFFFF1;
    // rom_array[31573] = 32'hFFFFFFF1;
    // rom_array[31574] = 32'hFFFFFFF1;
    // rom_array[31575] = 32'hFFFFFFF1;
    // rom_array[31576] = 32'hFFFFFFF1;
    // rom_array[31577] = 32'hFFFFFFF0;
    // rom_array[31578] = 32'hFFFFFFF0;
    // rom_array[31579] = 32'hFFFFFFF0;
    // rom_array[31580] = 32'hFFFFFFF0;
    // rom_array[31581] = 32'hFFFFFFF1;
    // rom_array[31582] = 32'hFFFFFFF1;
    // rom_array[31583] = 32'hFFFFFFF1;
    // rom_array[31584] = 32'hFFFFFFF1;
    // rom_array[31585] = 32'hFFFFFFF0;
    // rom_array[31586] = 32'hFFFFFFF0;
    // rom_array[31587] = 32'hFFFFFFF0;
    // rom_array[31588] = 32'hFFFFFFF0;
    // rom_array[31589] = 32'hFFFFFFF1;
    // rom_array[31590] = 32'hFFFFFFF1;
    // rom_array[31591] = 32'hFFFFFFF1;
    // rom_array[31592] = 32'hFFFFFFF1;
    // rom_array[31593] = 32'hFFFFFFF0;
    // rom_array[31594] = 32'hFFFFFFF0;
    // rom_array[31595] = 32'hFFFFFFF0;
    // rom_array[31596] = 32'hFFFFFFF0;
    // rom_array[31597] = 32'hFFFFFFF1;
    // rom_array[31598] = 32'hFFFFFFF1;
    // rom_array[31599] = 32'hFFFFFFF1;
    // rom_array[31600] = 32'hFFFFFFF1;
    // rom_array[31601] = 32'hFFFFFFF0;
    // rom_array[31602] = 32'hFFFFFFF0;
    // rom_array[31603] = 32'hFFFFFFF0;
    // rom_array[31604] = 32'hFFFFFFF0;
    // rom_array[31605] = 32'hFFFFFFF1;
    // rom_array[31606] = 32'hFFFFFFF1;
    // rom_array[31607] = 32'hFFFFFFF1;
    // rom_array[31608] = 32'hFFFFFFF1;
    // rom_array[31609] = 32'hFFFFFFF0;
    // rom_array[31610] = 32'hFFFFFFF0;
    // rom_array[31611] = 32'hFFFFFFF0;
    // rom_array[31612] = 32'hFFFFFFF0;
    // rom_array[31613] = 32'hFFFFFFF1;
    // rom_array[31614] = 32'hFFFFFFF1;
    // rom_array[31615] = 32'hFFFFFFF1;
    // rom_array[31616] = 32'hFFFFFFF1;
    // rom_array[31617] = 32'hFFFFFFF0;
    // rom_array[31618] = 32'hFFFFFFF0;
    // rom_array[31619] = 32'hFFFFFFF0;
    // rom_array[31620] = 32'hFFFFFFF0;
    // rom_array[31621] = 32'hFFFFFFF1;
    // rom_array[31622] = 32'hFFFFFFF1;
    // rom_array[31623] = 32'hFFFFFFF1;
    // rom_array[31624] = 32'hFFFFFFF1;
    // rom_array[31625] = 32'hFFFFFFF0;
    // rom_array[31626] = 32'hFFFFFFF0;
    // rom_array[31627] = 32'hFFFFFFF0;
    // rom_array[31628] = 32'hFFFFFFF0;
    // rom_array[31629] = 32'hFFFFFFF1;
    // rom_array[31630] = 32'hFFFFFFF1;
    // rom_array[31631] = 32'hFFFFFFF1;
    // rom_array[31632] = 32'hFFFFFFF1;
    // rom_array[31633] = 32'hFFFFFFF0;
    // rom_array[31634] = 32'hFFFFFFF0;
    // rom_array[31635] = 32'hFFFFFFF0;
    // rom_array[31636] = 32'hFFFFFFF0;
    // rom_array[31637] = 32'hFFFFFFF1;
    // rom_array[31638] = 32'hFFFFFFF1;
    // rom_array[31639] = 32'hFFFFFFF1;
    // rom_array[31640] = 32'hFFFFFFF1;
    // rom_array[31641] = 32'hFFFFFFF0;
    // rom_array[31642] = 32'hFFFFFFF0;
    // rom_array[31643] = 32'hFFFFFFF0;
    // rom_array[31644] = 32'hFFFFFFF0;
    // rom_array[31645] = 32'hFFFFFFF1;
    // rom_array[31646] = 32'hFFFFFFF1;
    // rom_array[31647] = 32'hFFFFFFF1;
    // rom_array[31648] = 32'hFFFFFFF1;
    // rom_array[31649] = 32'hFFFFFFF0;
    // rom_array[31650] = 32'hFFFFFFF0;
    // rom_array[31651] = 32'hFFFFFFF0;
    // rom_array[31652] = 32'hFFFFFFF0;
    // rom_array[31653] = 32'hFFFFFFF1;
    // rom_array[31654] = 32'hFFFFFFF1;
    // rom_array[31655] = 32'hFFFFFFF1;
    // rom_array[31656] = 32'hFFFFFFF1;
    // rom_array[31657] = 32'hFFFFFFF0;
    // rom_array[31658] = 32'hFFFFFFF0;
    // rom_array[31659] = 32'hFFFFFFF0;
    // rom_array[31660] = 32'hFFFFFFF0;
    // rom_array[31661] = 32'hFFFFFFF1;
    // rom_array[31662] = 32'hFFFFFFF1;
    // rom_array[31663] = 32'hFFFFFFF1;
    // rom_array[31664] = 32'hFFFFFFF1;
    // rom_array[31665] = 32'hFFFFFFF0;
    // rom_array[31666] = 32'hFFFFFFF0;
    // rom_array[31667] = 32'hFFFFFFF0;
    // rom_array[31668] = 32'hFFFFFFF0;
    // rom_array[31669] = 32'hFFFFFFF1;
    // rom_array[31670] = 32'hFFFFFFF1;
    // rom_array[31671] = 32'hFFFFFFF1;
    // rom_array[31672] = 32'hFFFFFFF1;
    // rom_array[31673] = 32'hFFFFFFF0;
    // rom_array[31674] = 32'hFFFFFFF0;
    // rom_array[31675] = 32'hFFFFFFF1;
    // rom_array[31676] = 32'hFFFFFFF1;
    // rom_array[31677] = 32'hFFFFFFF0;
    // rom_array[31678] = 32'hFFFFFFF0;
    // rom_array[31679] = 32'hFFFFFFF1;
    // rom_array[31680] = 32'hFFFFFFF1;
    // rom_array[31681] = 32'hFFFFFFF0;
    // rom_array[31682] = 32'hFFFFFFF0;
    // rom_array[31683] = 32'hFFFFFFF1;
    // rom_array[31684] = 32'hFFFFFFF1;
    // rom_array[31685] = 32'hFFFFFFF0;
    // rom_array[31686] = 32'hFFFFFFF0;
    // rom_array[31687] = 32'hFFFFFFF1;
    // rom_array[31688] = 32'hFFFFFFF1;
    // rom_array[31689] = 32'hFFFFFFF0;
    // rom_array[31690] = 32'hFFFFFFF0;
    // rom_array[31691] = 32'hFFFFFFF1;
    // rom_array[31692] = 32'hFFFFFFF1;
    // rom_array[31693] = 32'hFFFFFFF0;
    // rom_array[31694] = 32'hFFFFFFF0;
    // rom_array[31695] = 32'hFFFFFFF1;
    // rom_array[31696] = 32'hFFFFFFF1;
    // rom_array[31697] = 32'hFFFFFFF0;
    // rom_array[31698] = 32'hFFFFFFF0;
    // rom_array[31699] = 32'hFFFFFFF1;
    // rom_array[31700] = 32'hFFFFFFF1;
    // rom_array[31701] = 32'hFFFFFFF0;
    // rom_array[31702] = 32'hFFFFFFF0;
    // rom_array[31703] = 32'hFFFFFFF1;
    // rom_array[31704] = 32'hFFFFFFF1;
    // rom_array[31705] = 32'hFFFFFFF0;
    // rom_array[31706] = 32'hFFFFFFF0;
    // rom_array[31707] = 32'hFFFFFFF1;
    // rom_array[31708] = 32'hFFFFFFF1;
    // rom_array[31709] = 32'hFFFFFFF0;
    // rom_array[31710] = 32'hFFFFFFF0;
    // rom_array[31711] = 32'hFFFFFFF1;
    // rom_array[31712] = 32'hFFFFFFF1;
    // rom_array[31713] = 32'hFFFFFFF0;
    // rom_array[31714] = 32'hFFFFFFF0;
    // rom_array[31715] = 32'hFFFFFFF1;
    // rom_array[31716] = 32'hFFFFFFF1;
    // rom_array[31717] = 32'hFFFFFFF0;
    // rom_array[31718] = 32'hFFFFFFF0;
    // rom_array[31719] = 32'hFFFFFFF1;
    // rom_array[31720] = 32'hFFFFFFF1;
    // rom_array[31721] = 32'hFFFFFFF0;
    // rom_array[31722] = 32'hFFFFFFF0;
    // rom_array[31723] = 32'hFFFFFFF1;
    // rom_array[31724] = 32'hFFFFFFF1;
    // rom_array[31725] = 32'hFFFFFFF0;
    // rom_array[31726] = 32'hFFFFFFF0;
    // rom_array[31727] = 32'hFFFFFFF1;
    // rom_array[31728] = 32'hFFFFFFF1;
    // rom_array[31729] = 32'hFFFFFFF0;
    // rom_array[31730] = 32'hFFFFFFF0;
    // rom_array[31731] = 32'hFFFFFFF1;
    // rom_array[31732] = 32'hFFFFFFF1;
    // rom_array[31733] = 32'hFFFFFFF0;
    // rom_array[31734] = 32'hFFFFFFF0;
    // rom_array[31735] = 32'hFFFFFFF1;
    // rom_array[31736] = 32'hFFFFFFF1;
    // rom_array[31737] = 32'hFFFFFFF0;
    // rom_array[31738] = 32'hFFFFFFF0;
    // rom_array[31739] = 32'hFFFFFFF1;
    // rom_array[31740] = 32'hFFFFFFF1;
    // rom_array[31741] = 32'hFFFFFFF0;
    // rom_array[31742] = 32'hFFFFFFF0;
    // rom_array[31743] = 32'hFFFFFFF1;
    // rom_array[31744] = 32'hFFFFFFF1;
    // rom_array[31745] = 32'hFFFFFFF0;
    // rom_array[31746] = 32'hFFFFFFF0;
    // rom_array[31747] = 32'hFFFFFFF1;
    // rom_array[31748] = 32'hFFFFFFF1;
    // rom_array[31749] = 32'hFFFFFFF0;
    // rom_array[31750] = 32'hFFFFFFF0;
    // rom_array[31751] = 32'hFFFFFFF1;
    // rom_array[31752] = 32'hFFFFFFF1;
    // rom_array[31753] = 32'hFFFFFFF0;
    // rom_array[31754] = 32'hFFFFFFF0;
    // rom_array[31755] = 32'hFFFFFFF1;
    // rom_array[31756] = 32'hFFFFFFF1;
    // rom_array[31757] = 32'hFFFFFFF0;
    // rom_array[31758] = 32'hFFFFFFF0;
    // rom_array[31759] = 32'hFFFFFFF1;
    // rom_array[31760] = 32'hFFFFFFF1;
    // rom_array[31761] = 32'hFFFFFFF0;
    // rom_array[31762] = 32'hFFFFFFF0;
    // rom_array[31763] = 32'hFFFFFFF1;
    // rom_array[31764] = 32'hFFFFFFF1;
    // rom_array[31765] = 32'hFFFFFFF0;
    // rom_array[31766] = 32'hFFFFFFF0;
    // rom_array[31767] = 32'hFFFFFFF1;
    // rom_array[31768] = 32'hFFFFFFF1;
    // rom_array[31769] = 32'hFFFFFFF0;
    // rom_array[31770] = 32'hFFFFFFF0;
    // rom_array[31771] = 32'hFFFFFFF1;
    // rom_array[31772] = 32'hFFFFFFF1;
    // rom_array[31773] = 32'hFFFFFFF0;
    // rom_array[31774] = 32'hFFFFFFF0;
    // rom_array[31775] = 32'hFFFFFFF1;
    // rom_array[31776] = 32'hFFFFFFF1;
    // rom_array[31777] = 32'hFFFFFFF0;
    // rom_array[31778] = 32'hFFFFFFF0;
    // rom_array[31779] = 32'hFFFFFFF1;
    // rom_array[31780] = 32'hFFFFFFF1;
    // rom_array[31781] = 32'hFFFFFFF0;
    // rom_array[31782] = 32'hFFFFFFF0;
    // rom_array[31783] = 32'hFFFFFFF1;
    // rom_array[31784] = 32'hFFFFFFF1;
    // rom_array[31785] = 32'hFFFFFFF0;
    // rom_array[31786] = 32'hFFFFFFF0;
    // rom_array[31787] = 32'hFFFFFFF1;
    // rom_array[31788] = 32'hFFFFFFF1;
    // rom_array[31789] = 32'hFFFFFFF0;
    // rom_array[31790] = 32'hFFFFFFF0;
    // rom_array[31791] = 32'hFFFFFFF0;
    // rom_array[31792] = 32'hFFFFFFF0;
    // rom_array[31793] = 32'hFFFFFFF0;
    // rom_array[31794] = 32'hFFFFFFF0;
    // rom_array[31795] = 32'hFFFFFFF1;
    // rom_array[31796] = 32'hFFFFFFF1;
    // rom_array[31797] = 32'hFFFFFFF0;
    // rom_array[31798] = 32'hFFFFFFF0;
    // rom_array[31799] = 32'hFFFFFFF0;
    // rom_array[31800] = 32'hFFFFFFF0;
    // rom_array[31801] = 32'hFFFFFFF1;
    // rom_array[31802] = 32'hFFFFFFF1;
    // rom_array[31803] = 32'hFFFFFFF1;
    // rom_array[31804] = 32'hFFFFFFF1;
    // rom_array[31805] = 32'hFFFFFFF0;
    // rom_array[31806] = 32'hFFFFFFF0;
    // rom_array[31807] = 32'hFFFFFFF0;
    // rom_array[31808] = 32'hFFFFFFF0;
    // rom_array[31809] = 32'hFFFFFFF1;
    // rom_array[31810] = 32'hFFFFFFF1;
    // rom_array[31811] = 32'hFFFFFFF1;
    // rom_array[31812] = 32'hFFFFFFF1;
    // rom_array[31813] = 32'hFFFFFFF0;
    // rom_array[31814] = 32'hFFFFFFF0;
    // rom_array[31815] = 32'hFFFFFFF0;
    // rom_array[31816] = 32'hFFFFFFF0;
    // rom_array[31817] = 32'hFFFFFFF1;
    // rom_array[31818] = 32'hFFFFFFF1;
    // rom_array[31819] = 32'hFFFFFFF1;
    // rom_array[31820] = 32'hFFFFFFF1;
    // rom_array[31821] = 32'hFFFFFFF0;
    // rom_array[31822] = 32'hFFFFFFF0;
    // rom_array[31823] = 32'hFFFFFFF0;
    // rom_array[31824] = 32'hFFFFFFF0;
    // rom_array[31825] = 32'hFFFFFFF1;
    // rom_array[31826] = 32'hFFFFFFF1;
    // rom_array[31827] = 32'hFFFFFFF1;
    // rom_array[31828] = 32'hFFFFFFF1;
    // rom_array[31829] = 32'hFFFFFFF0;
    // rom_array[31830] = 32'hFFFFFFF0;
    // rom_array[31831] = 32'hFFFFFFF0;
    // rom_array[31832] = 32'hFFFFFFF0;
    // rom_array[31833] = 32'hFFFFFFF1;
    // rom_array[31834] = 32'hFFFFFFF1;
    // rom_array[31835] = 32'hFFFFFFF1;
    // rom_array[31836] = 32'hFFFFFFF1;
    // rom_array[31837] = 32'hFFFFFFF0;
    // rom_array[31838] = 32'hFFFFFFF0;
    // rom_array[31839] = 32'hFFFFFFF0;
    // rom_array[31840] = 32'hFFFFFFF0;
    // rom_array[31841] = 32'hFFFFFFF1;
    // rom_array[31842] = 32'hFFFFFFF1;
    // rom_array[31843] = 32'hFFFFFFF1;
    // rom_array[31844] = 32'hFFFFFFF1;
    // rom_array[31845] = 32'hFFFFFFF0;
    // rom_array[31846] = 32'hFFFFFFF0;
    // rom_array[31847] = 32'hFFFFFFF0;
    // rom_array[31848] = 32'hFFFFFFF0;
    // rom_array[31849] = 32'hFFFFFFF1;
    // rom_array[31850] = 32'hFFFFFFF1;
    // rom_array[31851] = 32'hFFFFFFF1;
    // rom_array[31852] = 32'hFFFFFFF1;
    // rom_array[31853] = 32'hFFFFFFF1;
    // rom_array[31854] = 32'hFFFFFFF1;
    // rom_array[31855] = 32'hFFFFFFF1;
    // rom_array[31856] = 32'hFFFFFFF1;
    // rom_array[31857] = 32'hFFFFFFF1;
    // rom_array[31858] = 32'hFFFFFFF1;
    // rom_array[31859] = 32'hFFFFFFF1;
    // rom_array[31860] = 32'hFFFFFFF1;
    // rom_array[31861] = 32'hFFFFFFF1;
    // rom_array[31862] = 32'hFFFFFFF1;
    // rom_array[31863] = 32'hFFFFFFF1;
    // rom_array[31864] = 32'hFFFFFFF1;
    // rom_array[31865] = 32'hFFFFFFF1;
    // rom_array[31866] = 32'hFFFFFFF1;
    // rom_array[31867] = 32'hFFFFFFF1;
    // rom_array[31868] = 32'hFFFFFFF1;
    // rom_array[31869] = 32'hFFFFFFF1;
    // rom_array[31870] = 32'hFFFFFFF1;
    // rom_array[31871] = 32'hFFFFFFF1;
    // rom_array[31872] = 32'hFFFFFFF1;
    // rom_array[31873] = 32'hFFFFFFF1;
    // rom_array[31874] = 32'hFFFFFFF1;
    // rom_array[31875] = 32'hFFFFFFF1;
    // rom_array[31876] = 32'hFFFFFFF1;
    // rom_array[31877] = 32'hFFFFFFF1;
    // rom_array[31878] = 32'hFFFFFFF1;
    // rom_array[31879] = 32'hFFFFFFF1;
    // rom_array[31880] = 32'hFFFFFFF1;
    // rom_array[31881] = 32'hFFFFFFF1;
    // rom_array[31882] = 32'hFFFFFFF1;
    // rom_array[31883] = 32'hFFFFFFF1;
    // rom_array[31884] = 32'hFFFFFFF1;
    // rom_array[31885] = 32'hFFFFFFF1;
    // rom_array[31886] = 32'hFFFFFFF1;
    // rom_array[31887] = 32'hFFFFFFF1;
    // rom_array[31888] = 32'hFFFFFFF1;
    // rom_array[31889] = 32'hFFFFFFF1;
    // rom_array[31890] = 32'hFFFFFFF1;
    // rom_array[31891] = 32'hFFFFFFF1;
    // rom_array[31892] = 32'hFFFFFFF1;
    // rom_array[31893] = 32'hFFFFFFF1;
    // rom_array[31894] = 32'hFFFFFFF1;
    // rom_array[31895] = 32'hFFFFFFF1;
    // rom_array[31896] = 32'hFFFFFFF1;
    // rom_array[31897] = 32'hFFFFFFF1;
    // rom_array[31898] = 32'hFFFFFFF1;
    // rom_array[31899] = 32'hFFFFFFF1;
    // rom_array[31900] = 32'hFFFFFFF1;
    // rom_array[31901] = 32'hFFFFFFF0;
    // rom_array[31902] = 32'hFFFFFFF0;
    // rom_array[31903] = 32'hFFFFFFF0;
    // rom_array[31904] = 32'hFFFFFFF0;
    // rom_array[31905] = 32'hFFFFFFF1;
    // rom_array[31906] = 32'hFFFFFFF1;
    // rom_array[31907] = 32'hFFFFFFF1;
    // rom_array[31908] = 32'hFFFFFFF1;
    // rom_array[31909] = 32'hFFFFFFF0;
    // rom_array[31910] = 32'hFFFFFFF0;
    // rom_array[31911] = 32'hFFFFFFF0;
    // rom_array[31912] = 32'hFFFFFFF0;
    // rom_array[31913] = 32'hFFFFFFF1;
    // rom_array[31914] = 32'hFFFFFFF1;
    // rom_array[31915] = 32'hFFFFFFF1;
    // rom_array[31916] = 32'hFFFFFFF1;
    // rom_array[31917] = 32'hFFFFFFF1;
    // rom_array[31918] = 32'hFFFFFFF1;
    // rom_array[31919] = 32'hFFFFFFF1;
    // rom_array[31920] = 32'hFFFFFFF1;
    // rom_array[31921] = 32'hFFFFFFF1;
    // rom_array[31922] = 32'hFFFFFFF1;
    // rom_array[31923] = 32'hFFFFFFF1;
    // rom_array[31924] = 32'hFFFFFFF1;
    // rom_array[31925] = 32'hFFFFFFF1;
    // rom_array[31926] = 32'hFFFFFFF1;
    // rom_array[31927] = 32'hFFFFFFF1;
    // rom_array[31928] = 32'hFFFFFFF1;
    // rom_array[31929] = 32'hFFFFFFF1;
    // rom_array[31930] = 32'hFFFFFFF1;
    // rom_array[31931] = 32'hFFFFFFF1;
    // rom_array[31932] = 32'hFFFFFFF1;
    // rom_array[31933] = 32'hFFFFFFF0;
    // rom_array[31934] = 32'hFFFFFFF0;
    // rom_array[31935] = 32'hFFFFFFF0;
    // rom_array[31936] = 32'hFFFFFFF0;
    // rom_array[31937] = 32'hFFFFFFF1;
    // rom_array[31938] = 32'hFFFFFFF1;
    // rom_array[31939] = 32'hFFFFFFF1;
    // rom_array[31940] = 32'hFFFFFFF1;
    // rom_array[31941] = 32'hFFFFFFF0;
    // rom_array[31942] = 32'hFFFFFFF0;
    // rom_array[31943] = 32'hFFFFFFF0;
    // rom_array[31944] = 32'hFFFFFFF0;
    // rom_array[31945] = 32'hFFFFFFF1;
    // rom_array[31946] = 32'hFFFFFFF1;
    // rom_array[31947] = 32'hFFFFFFF1;
    // rom_array[31948] = 32'hFFFFFFF1;
    // rom_array[31949] = 32'hFFFFFFF0;
    // rom_array[31950] = 32'hFFFFFFF0;
    // rom_array[31951] = 32'hFFFFFFF0;
    // rom_array[31952] = 32'hFFFFFFF0;
    // rom_array[31953] = 32'hFFFFFFF1;
    // rom_array[31954] = 32'hFFFFFFF1;
    // rom_array[31955] = 32'hFFFFFFF1;
    // rom_array[31956] = 32'hFFFFFFF1;
    // rom_array[31957] = 32'hFFFFFFF0;
    // rom_array[31958] = 32'hFFFFFFF0;
    // rom_array[31959] = 32'hFFFFFFF0;
    // rom_array[31960] = 32'hFFFFFFF0;
    // rom_array[31961] = 32'hFFFFFFF1;
    // rom_array[31962] = 32'hFFFFFFF1;
    // rom_array[31963] = 32'hFFFFFFF1;
    // rom_array[31964] = 32'hFFFFFFF1;
    // rom_array[31965] = 32'hFFFFFFF0;
    // rom_array[31966] = 32'hFFFFFFF0;
    // rom_array[31967] = 32'hFFFFFFF0;
    // rom_array[31968] = 32'hFFFFFFF0;
    // rom_array[31969] = 32'hFFFFFFF1;
    // rom_array[31970] = 32'hFFFFFFF1;
    // rom_array[31971] = 32'hFFFFFFF1;
    // rom_array[31972] = 32'hFFFFFFF1;
    // rom_array[31973] = 32'hFFFFFFF0;
    // rom_array[31974] = 32'hFFFFFFF0;
    // rom_array[31975] = 32'hFFFFFFF0;
    // rom_array[31976] = 32'hFFFFFFF0;
    // rom_array[31977] = 32'hFFFFFFF1;
    // rom_array[31978] = 32'hFFFFFFF1;
    // rom_array[31979] = 32'hFFFFFFF1;
    // rom_array[31980] = 32'hFFFFFFF1;
    // rom_array[31981] = 32'hFFFFFFF0;
    // rom_array[31982] = 32'hFFFFFFF0;
    // rom_array[31983] = 32'hFFFFFFF0;
    // rom_array[31984] = 32'hFFFFFFF0;
    // rom_array[31985] = 32'hFFFFFFF1;
    // rom_array[31986] = 32'hFFFFFFF1;
    // rom_array[31987] = 32'hFFFFFFF1;
    // rom_array[31988] = 32'hFFFFFFF1;
    // rom_array[31989] = 32'hFFFFFFF0;
    // rom_array[31990] = 32'hFFFFFFF0;
    // rom_array[31991] = 32'hFFFFFFF0;
    // rom_array[31992] = 32'hFFFFFFF0;
    // rom_array[31993] = 32'hFFFFFFF1;
    // rom_array[31994] = 32'hFFFFFFF1;
    // rom_array[31995] = 32'hFFFFFFF1;
    // rom_array[31996] = 32'hFFFFFFF1;
    // rom_array[31997] = 32'hFFFFFFF0;
    // rom_array[31998] = 32'hFFFFFFF0;
    // rom_array[31999] = 32'hFFFFFFF0;
    // rom_array[32000] = 32'hFFFFFFF0;
    // rom_array[32001] = 32'hFFFFFFF1;
    // rom_array[32002] = 32'hFFFFFFF1;
    // rom_array[32003] = 32'hFFFFFFF1;
    // rom_array[32004] = 32'hFFFFFFF1;
    // rom_array[32005] = 32'hFFFFFFF0;
    // rom_array[32006] = 32'hFFFFFFF0;
    // rom_array[32007] = 32'hFFFFFFF0;
    // rom_array[32008] = 32'hFFFFFFF0;
    // rom_array[32009] = 32'hFFFFFFF1;
    // rom_array[32010] = 32'hFFFFFFF1;
    // rom_array[32011] = 32'hFFFFFFF1;
    // rom_array[32012] = 32'hFFFFFFF1;
    // rom_array[32013] = 32'hFFFFFFF0;
    // rom_array[32014] = 32'hFFFFFFF0;
    // rom_array[32015] = 32'hFFFFFFF0;
    // rom_array[32016] = 32'hFFFFFFF0;
    // rom_array[32017] = 32'hFFFFFFF1;
    // rom_array[32018] = 32'hFFFFFFF1;
    // rom_array[32019] = 32'hFFFFFFF1;
    // rom_array[32020] = 32'hFFFFFFF1;
    // rom_array[32021] = 32'hFFFFFFF0;
    // rom_array[32022] = 32'hFFFFFFF0;
    // rom_array[32023] = 32'hFFFFFFF0;
    // rom_array[32024] = 32'hFFFFFFF0;
    // rom_array[32025] = 32'hFFFFFFF1;
    // rom_array[32026] = 32'hFFFFFFF1;
    // rom_array[32027] = 32'hFFFFFFF1;
    // rom_array[32028] = 32'hFFFFFFF1;
    // rom_array[32029] = 32'hFFFFFFF1;
    // rom_array[32030] = 32'hFFFFFFF1;
    // rom_array[32031] = 32'hFFFFFFF1;
    // rom_array[32032] = 32'hFFFFFFF1;
    // rom_array[32033] = 32'hFFFFFFF1;
    // rom_array[32034] = 32'hFFFFFFF1;
    // rom_array[32035] = 32'hFFFFFFF1;
    // rom_array[32036] = 32'hFFFFFFF1;
    // rom_array[32037] = 32'hFFFFFFF1;
    // rom_array[32038] = 32'hFFFFFFF1;
    // rom_array[32039] = 32'hFFFFFFF1;
    // rom_array[32040] = 32'hFFFFFFF1;
    // rom_array[32041] = 32'hFFFFFFF1;
    // rom_array[32042] = 32'hFFFFFFF1;
    // rom_array[32043] = 32'hFFFFFFF1;
    // rom_array[32044] = 32'hFFFFFFF1;
    // rom_array[32045] = 32'hFFFFFFF1;
    // rom_array[32046] = 32'hFFFFFFF1;
    // rom_array[32047] = 32'hFFFFFFF1;
    // rom_array[32048] = 32'hFFFFFFF1;
    // rom_array[32049] = 32'hFFFFFFF1;
    // rom_array[32050] = 32'hFFFFFFF1;
    // rom_array[32051] = 32'hFFFFFFF1;
    // rom_array[32052] = 32'hFFFFFFF1;
    // rom_array[32053] = 32'hFFFFFFF1;
    // rom_array[32054] = 32'hFFFFFFF1;
    // rom_array[32055] = 32'hFFFFFFF1;
    // rom_array[32056] = 32'hFFFFFFF1;
    // rom_array[32057] = 32'hFFFFFFF1;
    // rom_array[32058] = 32'hFFFFFFF1;
    // rom_array[32059] = 32'hFFFFFFF1;
    // rom_array[32060] = 32'hFFFFFFF1;
    // rom_array[32061] = 32'hFFFFFFF1;
    // rom_array[32062] = 32'hFFFFFFF1;
    // rom_array[32063] = 32'hFFFFFFF1;
    // rom_array[32064] = 32'hFFFFFFF1;
    // rom_array[32065] = 32'hFFFFFFF1;
    // rom_array[32066] = 32'hFFFFFFF1;
    // rom_array[32067] = 32'hFFFFFFF1;
    // rom_array[32068] = 32'hFFFFFFF1;
    // rom_array[32069] = 32'hFFFFFFF1;
    // rom_array[32070] = 32'hFFFFFFF1;
    // rom_array[32071] = 32'hFFFFFFF1;
    // rom_array[32072] = 32'hFFFFFFF1;
    // rom_array[32073] = 32'hFFFFFFF1;
    // rom_array[32074] = 32'hFFFFFFF1;
    // rom_array[32075] = 32'hFFFFFFF1;
    // rom_array[32076] = 32'hFFFFFFF1;
    // rom_array[32077] = 32'hFFFFFFF0;
    // rom_array[32078] = 32'hFFFFFFF0;
    // rom_array[32079] = 32'hFFFFFFF0;
    // rom_array[32080] = 32'hFFFFFFF0;
    // rom_array[32081] = 32'hFFFFFFF1;
    // rom_array[32082] = 32'hFFFFFFF1;
    // rom_array[32083] = 32'hFFFFFFF1;
    // rom_array[32084] = 32'hFFFFFFF1;
    // rom_array[32085] = 32'hFFFFFFF0;
    // rom_array[32086] = 32'hFFFFFFF0;
    // rom_array[32087] = 32'hFFFFFFF0;
    // rom_array[32088] = 32'hFFFFFFF0;
    // rom_array[32089] = 32'hFFFFFFF0;
    // rom_array[32090] = 32'hFFFFFFF0;
    // rom_array[32091] = 32'hFFFFFFF0;
    // rom_array[32092] = 32'hFFFFFFF0;
    // rom_array[32093] = 32'hFFFFFFF0;
    // rom_array[32094] = 32'hFFFFFFF0;
    // rom_array[32095] = 32'hFFFFFFF1;
    // rom_array[32096] = 32'hFFFFFFF1;
    // rom_array[32097] = 32'hFFFFFFF0;
    // rom_array[32098] = 32'hFFFFFFF0;
    // rom_array[32099] = 32'hFFFFFFF0;
    // rom_array[32100] = 32'hFFFFFFF0;
    // rom_array[32101] = 32'hFFFFFFF0;
    // rom_array[32102] = 32'hFFFFFFF0;
    // rom_array[32103] = 32'hFFFFFFF1;
    // rom_array[32104] = 32'hFFFFFFF1;
    // rom_array[32105] = 32'hFFFFFFF0;
    // rom_array[32106] = 32'hFFFFFFF0;
    // rom_array[32107] = 32'hFFFFFFF0;
    // rom_array[32108] = 32'hFFFFFFF0;
    // rom_array[32109] = 32'hFFFFFFF1;
    // rom_array[32110] = 32'hFFFFFFF1;
    // rom_array[32111] = 32'hFFFFFFF1;
    // rom_array[32112] = 32'hFFFFFFF1;
    // rom_array[32113] = 32'hFFFFFFF0;
    // rom_array[32114] = 32'hFFFFFFF0;
    // rom_array[32115] = 32'hFFFFFFF0;
    // rom_array[32116] = 32'hFFFFFFF0;
    // rom_array[32117] = 32'hFFFFFFF1;
    // rom_array[32118] = 32'hFFFFFFF1;
    // rom_array[32119] = 32'hFFFFFFF1;
    // rom_array[32120] = 32'hFFFFFFF1;
    // rom_array[32121] = 32'hFFFFFFF0;
    // rom_array[32122] = 32'hFFFFFFF0;
    // rom_array[32123] = 32'hFFFFFFF1;
    // rom_array[32124] = 32'hFFFFFFF1;
    // rom_array[32125] = 32'hFFFFFFF0;
    // rom_array[32126] = 32'hFFFFFFF0;
    // rom_array[32127] = 32'hFFFFFFF1;
    // rom_array[32128] = 32'hFFFFFFF1;
    // rom_array[32129] = 32'hFFFFFFF0;
    // rom_array[32130] = 32'hFFFFFFF0;
    // rom_array[32131] = 32'hFFFFFFF1;
    // rom_array[32132] = 32'hFFFFFFF1;
    // rom_array[32133] = 32'hFFFFFFF0;
    // rom_array[32134] = 32'hFFFFFFF0;
    // rom_array[32135] = 32'hFFFFFFF1;
    // rom_array[32136] = 32'hFFFFFFF1;
    // rom_array[32137] = 32'hFFFFFFF0;
    // rom_array[32138] = 32'hFFFFFFF0;
    // rom_array[32139] = 32'hFFFFFFF0;
    // rom_array[32140] = 32'hFFFFFFF0;
    // rom_array[32141] = 32'hFFFFFFF1;
    // rom_array[32142] = 32'hFFFFFFF1;
    // rom_array[32143] = 32'hFFFFFFF1;
    // rom_array[32144] = 32'hFFFFFFF1;
    // rom_array[32145] = 32'hFFFFFFF0;
    // rom_array[32146] = 32'hFFFFFFF0;
    // rom_array[32147] = 32'hFFFFFFF0;
    // rom_array[32148] = 32'hFFFFFFF0;
    // rom_array[32149] = 32'hFFFFFFF1;
    // rom_array[32150] = 32'hFFFFFFF1;
    // rom_array[32151] = 32'hFFFFFFF1;
    // rom_array[32152] = 32'hFFFFFFF1;
    // rom_array[32153] = 32'hFFFFFFF0;
    // rom_array[32154] = 32'hFFFFFFF0;
    // rom_array[32155] = 32'hFFFFFFF0;
    // rom_array[32156] = 32'hFFFFFFF0;
    // rom_array[32157] = 32'hFFFFFFF1;
    // rom_array[32158] = 32'hFFFFFFF1;
    // rom_array[32159] = 32'hFFFFFFF1;
    // rom_array[32160] = 32'hFFFFFFF1;
    // rom_array[32161] = 32'hFFFFFFF0;
    // rom_array[32162] = 32'hFFFFFFF0;
    // rom_array[32163] = 32'hFFFFFFF0;
    // rom_array[32164] = 32'hFFFFFFF0;
    // rom_array[32165] = 32'hFFFFFFF1;
    // rom_array[32166] = 32'hFFFFFFF1;
    // rom_array[32167] = 32'hFFFFFFF1;
    // rom_array[32168] = 32'hFFFFFFF1;
    // rom_array[32169] = 32'hFFFFFFF0;
    // rom_array[32170] = 32'hFFFFFFF0;
    // rom_array[32171] = 32'hFFFFFFF0;
    // rom_array[32172] = 32'hFFFFFFF0;
    // rom_array[32173] = 32'hFFFFFFF1;
    // rom_array[32174] = 32'hFFFFFFF1;
    // rom_array[32175] = 32'hFFFFFFF1;
    // rom_array[32176] = 32'hFFFFFFF1;
    // rom_array[32177] = 32'hFFFFFFF0;
    // rom_array[32178] = 32'hFFFFFFF0;
    // rom_array[32179] = 32'hFFFFFFF0;
    // rom_array[32180] = 32'hFFFFFFF0;
    // rom_array[32181] = 32'hFFFFFFF1;
    // rom_array[32182] = 32'hFFFFFFF1;
    // rom_array[32183] = 32'hFFFFFFF1;
    // rom_array[32184] = 32'hFFFFFFF1;
    // rom_array[32185] = 32'hFFFFFFF1;
    // rom_array[32186] = 32'hFFFFFFF1;
    // rom_array[32187] = 32'hFFFFFFF0;
    // rom_array[32188] = 32'hFFFFFFF0;
    // rom_array[32189] = 32'hFFFFFFF1;
    // rom_array[32190] = 32'hFFFFFFF1;
    // rom_array[32191] = 32'hFFFFFFF1;
    // rom_array[32192] = 32'hFFFFFFF1;
    // rom_array[32193] = 32'hFFFFFFF1;
    // rom_array[32194] = 32'hFFFFFFF1;
    // rom_array[32195] = 32'hFFFFFFF0;
    // rom_array[32196] = 32'hFFFFFFF0;
    // rom_array[32197] = 32'hFFFFFFF1;
    // rom_array[32198] = 32'hFFFFFFF1;
    // rom_array[32199] = 32'hFFFFFFF1;
    // rom_array[32200] = 32'hFFFFFFF1;
    // rom_array[32201] = 32'hFFFFFFF0;
    // rom_array[32202] = 32'hFFFFFFF0;
    // rom_array[32203] = 32'hFFFFFFF1;
    // rom_array[32204] = 32'hFFFFFFF1;
    // rom_array[32205] = 32'hFFFFFFF0;
    // rom_array[32206] = 32'hFFFFFFF0;
    // rom_array[32207] = 32'hFFFFFFF1;
    // rom_array[32208] = 32'hFFFFFFF1;
    // rom_array[32209] = 32'hFFFFFFF0;
    // rom_array[32210] = 32'hFFFFFFF0;
    // rom_array[32211] = 32'hFFFFFFF1;
    // rom_array[32212] = 32'hFFFFFFF1;
    // rom_array[32213] = 32'hFFFFFFF0;
    // rom_array[32214] = 32'hFFFFFFF0;
    // rom_array[32215] = 32'hFFFFFFF1;
    // rom_array[32216] = 32'hFFFFFFF1;
    // rom_array[32217] = 32'hFFFFFFF0;
    // rom_array[32218] = 32'hFFFFFFF0;
    // rom_array[32219] = 32'hFFFFFFF1;
    // rom_array[32220] = 32'hFFFFFFF1;
    // rom_array[32221] = 32'hFFFFFFF0;
    // rom_array[32222] = 32'hFFFFFFF0;
    // rom_array[32223] = 32'hFFFFFFF1;
    // rom_array[32224] = 32'hFFFFFFF1;
    // rom_array[32225] = 32'hFFFFFFF0;
    // rom_array[32226] = 32'hFFFFFFF0;
    // rom_array[32227] = 32'hFFFFFFF1;
    // rom_array[32228] = 32'hFFFFFFF1;
    // rom_array[32229] = 32'hFFFFFFF0;
    // rom_array[32230] = 32'hFFFFFFF0;
    // rom_array[32231] = 32'hFFFFFFF1;
    // rom_array[32232] = 32'hFFFFFFF1;
    // rom_array[32233] = 32'hFFFFFFF1;
    // rom_array[32234] = 32'hFFFFFFF1;
    // rom_array[32235] = 32'hFFFFFFF1;
    // rom_array[32236] = 32'hFFFFFFF1;
    // rom_array[32237] = 32'hFFFFFFF1;
    // rom_array[32238] = 32'hFFFFFFF1;
    // rom_array[32239] = 32'hFFFFFFF1;
    // rom_array[32240] = 32'hFFFFFFF1;
    // rom_array[32241] = 32'hFFFFFFF1;
    // rom_array[32242] = 32'hFFFFFFF1;
    // rom_array[32243] = 32'hFFFFFFF1;
    // rom_array[32244] = 32'hFFFFFFF1;
    // rom_array[32245] = 32'hFFFFFFF1;
    // rom_array[32246] = 32'hFFFFFFF1;
    // rom_array[32247] = 32'hFFFFFFF1;
    // rom_array[32248] = 32'hFFFFFFF1;
    // rom_array[32249] = 32'hFFFFFFF1;
    // rom_array[32250] = 32'hFFFFFFF1;
    // rom_array[32251] = 32'hFFFFFFF1;
    // rom_array[32252] = 32'hFFFFFFF1;
    // rom_array[32253] = 32'hFFFFFFF1;
    // rom_array[32254] = 32'hFFFFFFF1;
    // rom_array[32255] = 32'hFFFFFFF1;
    // rom_array[32256] = 32'hFFFFFFF1;
    // rom_array[32257] = 32'hFFFFFFF1;
    // rom_array[32258] = 32'hFFFFFFF1;
    // rom_array[32259] = 32'hFFFFFFF1;
    // rom_array[32260] = 32'hFFFFFFF1;
    // rom_array[32261] = 32'hFFFFFFF1;
    // rom_array[32262] = 32'hFFFFFFF1;
    // rom_array[32263] = 32'hFFFFFFF1;
    // rom_array[32264] = 32'hFFFFFFF1;
    // rom_array[32265] = 32'hFFFFFFF1;
    // rom_array[32266] = 32'hFFFFFFF1;
    // rom_array[32267] = 32'hFFFFFFF1;
    // rom_array[32268] = 32'hFFFFFFF1;
    // rom_array[32269] = 32'hFFFFFFF1;
    // rom_array[32270] = 32'hFFFFFFF1;
    // rom_array[32271] = 32'hFFFFFFF1;
    // rom_array[32272] = 32'hFFFFFFF1;
    // rom_array[32273] = 32'hFFFFFFF1;
    // rom_array[32274] = 32'hFFFFFFF1;
    // rom_array[32275] = 32'hFFFFFFF1;
    // rom_array[32276] = 32'hFFFFFFF1;
    // rom_array[32277] = 32'hFFFFFFF1;
    // rom_array[32278] = 32'hFFFFFFF1;
    // rom_array[32279] = 32'hFFFFFFF1;
    // rom_array[32280] = 32'hFFFFFFF1;
    // rom_array[32281] = 32'hFFFFFFF0;
    // rom_array[32282] = 32'hFFFFFFF0;
    // rom_array[32283] = 32'hFFFFFFF1;
    // rom_array[32284] = 32'hFFFFFFF1;
    // rom_array[32285] = 32'hFFFFFFF0;
    // rom_array[32286] = 32'hFFFFFFF0;
    // rom_array[32287] = 32'hFFFFFFF1;
    // rom_array[32288] = 32'hFFFFFFF1;
    // rom_array[32289] = 32'hFFFFFFF0;
    // rom_array[32290] = 32'hFFFFFFF0;
    // rom_array[32291] = 32'hFFFFFFF1;
    // rom_array[32292] = 32'hFFFFFFF1;
    // rom_array[32293] = 32'hFFFFFFF0;
    // rom_array[32294] = 32'hFFFFFFF0;
    // rom_array[32295] = 32'hFFFFFFF1;
    // rom_array[32296] = 32'hFFFFFFF1;
    // rom_array[32297] = 32'hFFFFFFF1;
    // rom_array[32298] = 32'hFFFFFFF1;
    // rom_array[32299] = 32'hFFFFFFF1;
    // rom_array[32300] = 32'hFFFFFFF1;
    // rom_array[32301] = 32'hFFFFFFF1;
    // rom_array[32302] = 32'hFFFFFFF1;
    // rom_array[32303] = 32'hFFFFFFF1;
    // rom_array[32304] = 32'hFFFFFFF1;
    // rom_array[32305] = 32'hFFFFFFF1;
    // rom_array[32306] = 32'hFFFFFFF1;
    // rom_array[32307] = 32'hFFFFFFF1;
    // rom_array[32308] = 32'hFFFFFFF1;
    // rom_array[32309] = 32'hFFFFFFF1;
    // rom_array[32310] = 32'hFFFFFFF1;
    // rom_array[32311] = 32'hFFFFFFF1;
    // rom_array[32312] = 32'hFFFFFFF1;
    // rom_array[32313] = 32'hFFFFFFF0;
    // rom_array[32314] = 32'hFFFFFFF0;
    // rom_array[32315] = 32'hFFFFFFF1;
    // rom_array[32316] = 32'hFFFFFFF1;
    // rom_array[32317] = 32'hFFFFFFF0;
    // rom_array[32318] = 32'hFFFFFFF0;
    // rom_array[32319] = 32'hFFFFFFF1;
    // rom_array[32320] = 32'hFFFFFFF1;
    // rom_array[32321] = 32'hFFFFFFF0;
    // rom_array[32322] = 32'hFFFFFFF0;
    // rom_array[32323] = 32'hFFFFFFF1;
    // rom_array[32324] = 32'hFFFFFFF1;
    // rom_array[32325] = 32'hFFFFFFF0;
    // rom_array[32326] = 32'hFFFFFFF0;
    // rom_array[32327] = 32'hFFFFFFF1;
    // rom_array[32328] = 32'hFFFFFFF1;
    // rom_array[32329] = 32'hFFFFFFF1;
    // rom_array[32330] = 32'hFFFFFFF1;
    // rom_array[32331] = 32'hFFFFFFF1;
    // rom_array[32332] = 32'hFFFFFFF1;
    // rom_array[32333] = 32'hFFFFFFF1;
    // rom_array[32334] = 32'hFFFFFFF1;
    // rom_array[32335] = 32'hFFFFFFF1;
    // rom_array[32336] = 32'hFFFFFFF1;
    // rom_array[32337] = 32'hFFFFFFF1;
    // rom_array[32338] = 32'hFFFFFFF1;
    // rom_array[32339] = 32'hFFFFFFF1;
    // rom_array[32340] = 32'hFFFFFFF1;
    // rom_array[32341] = 32'hFFFFFFF1;
    // rom_array[32342] = 32'hFFFFFFF1;
    // rom_array[32343] = 32'hFFFFFFF1;
    // rom_array[32344] = 32'hFFFFFFF1;
    // rom_array[32345] = 32'hFFFFFFF0;
    // rom_array[32346] = 32'hFFFFFFF0;
    // rom_array[32347] = 32'hFFFFFFF1;
    // rom_array[32348] = 32'hFFFFFFF1;
    // rom_array[32349] = 32'hFFFFFFF0;
    // rom_array[32350] = 32'hFFFFFFF0;
    // rom_array[32351] = 32'hFFFFFFF1;
    // rom_array[32352] = 32'hFFFFFFF1;
    // rom_array[32353] = 32'hFFFFFFF0;
    // rom_array[32354] = 32'hFFFFFFF0;
    // rom_array[32355] = 32'hFFFFFFF1;
    // rom_array[32356] = 32'hFFFFFFF1;
    // rom_array[32357] = 32'hFFFFFFF0;
    // rom_array[32358] = 32'hFFFFFFF0;
    // rom_array[32359] = 32'hFFFFFFF1;
    // rom_array[32360] = 32'hFFFFFFF1;
    // rom_array[32361] = 32'hFFFFFFF0;
    // rom_array[32362] = 32'hFFFFFFF0;
    // rom_array[32363] = 32'hFFFFFFF1;
    // rom_array[32364] = 32'hFFFFFFF1;
    // rom_array[32365] = 32'hFFFFFFF0;
    // rom_array[32366] = 32'hFFFFFFF0;
    // rom_array[32367] = 32'hFFFFFFF1;
    // rom_array[32368] = 32'hFFFFFFF1;
    // rom_array[32369] = 32'hFFFFFFF0;
    // rom_array[32370] = 32'hFFFFFFF0;
    // rom_array[32371] = 32'hFFFFFFF1;
    // rom_array[32372] = 32'hFFFFFFF1;
    // rom_array[32373] = 32'hFFFFFFF0;
    // rom_array[32374] = 32'hFFFFFFF0;
    // rom_array[32375] = 32'hFFFFFFF1;
    // rom_array[32376] = 32'hFFFFFFF1;
    // rom_array[32377] = 32'hFFFFFFF0;
    // rom_array[32378] = 32'hFFFFFFF0;
    // rom_array[32379] = 32'hFFFFFFF0;
    // rom_array[32380] = 32'hFFFFFFF0;
    // rom_array[32381] = 32'hFFFFFFF1;
    // rom_array[32382] = 32'hFFFFFFF1;
    // rom_array[32383] = 32'hFFFFFFF1;
    // rom_array[32384] = 32'hFFFFFFF1;
    // rom_array[32385] = 32'hFFFFFFF0;
    // rom_array[32386] = 32'hFFFFFFF0;
    // rom_array[32387] = 32'hFFFFFFF0;
    // rom_array[32388] = 32'hFFFFFFF0;
    // rom_array[32389] = 32'hFFFFFFF1;
    // rom_array[32390] = 32'hFFFFFFF1;
    // rom_array[32391] = 32'hFFFFFFF1;
    // rom_array[32392] = 32'hFFFFFFF1;
    // rom_array[32393] = 32'hFFFFFFF0;
    // rom_array[32394] = 32'hFFFFFFF0;
    // rom_array[32395] = 32'hFFFFFFF0;
    // rom_array[32396] = 32'hFFFFFFF0;
    // rom_array[32397] = 32'hFFFFFFF1;
    // rom_array[32398] = 32'hFFFFFFF1;
    // rom_array[32399] = 32'hFFFFFFF1;
    // rom_array[32400] = 32'hFFFFFFF1;
    // rom_array[32401] = 32'hFFFFFFF0;
    // rom_array[32402] = 32'hFFFFFFF0;
    // rom_array[32403] = 32'hFFFFFFF0;
    // rom_array[32404] = 32'hFFFFFFF0;
    // rom_array[32405] = 32'hFFFFFFF1;
    // rom_array[32406] = 32'hFFFFFFF1;
    // rom_array[32407] = 32'hFFFFFFF1;
    // rom_array[32408] = 32'hFFFFFFF1;
    // rom_array[32409] = 32'hFFFFFFF0;
    // rom_array[32410] = 32'hFFFFFFF0;
    // rom_array[32411] = 32'hFFFFFFF0;
    // rom_array[32412] = 32'hFFFFFFF0;
    // rom_array[32413] = 32'hFFFFFFF1;
    // rom_array[32414] = 32'hFFFFFFF1;
    // rom_array[32415] = 32'hFFFFFFF1;
    // rom_array[32416] = 32'hFFFFFFF1;
    // rom_array[32417] = 32'hFFFFFFF0;
    // rom_array[32418] = 32'hFFFFFFF0;
    // rom_array[32419] = 32'hFFFFFFF0;
    // rom_array[32420] = 32'hFFFFFFF0;
    // rom_array[32421] = 32'hFFFFFFF1;
    // rom_array[32422] = 32'hFFFFFFF1;
    // rom_array[32423] = 32'hFFFFFFF1;
    // rom_array[32424] = 32'hFFFFFFF1;
    // rom_array[32425] = 32'hFFFFFFF0;
    // rom_array[32426] = 32'hFFFFFFF0;
    // rom_array[32427] = 32'hFFFFFFF0;
    // rom_array[32428] = 32'hFFFFFFF0;
    // rom_array[32429] = 32'hFFFFFFF1;
    // rom_array[32430] = 32'hFFFFFFF1;
    // rom_array[32431] = 32'hFFFFFFF1;
    // rom_array[32432] = 32'hFFFFFFF1;
    // rom_array[32433] = 32'hFFFFFFF0;
    // rom_array[32434] = 32'hFFFFFFF0;
    // rom_array[32435] = 32'hFFFFFFF0;
    // rom_array[32436] = 32'hFFFFFFF0;
    // rom_array[32437] = 32'hFFFFFFF1;
    // rom_array[32438] = 32'hFFFFFFF1;
    // rom_array[32439] = 32'hFFFFFFF1;
    // rom_array[32440] = 32'hFFFFFFF1;
    // rom_array[32441] = 32'hFFFFFFF0;
    // rom_array[32442] = 32'hFFFFFFF0;
    // rom_array[32443] = 32'hFFFFFFF0;
    // rom_array[32444] = 32'hFFFFFFF0;
    // rom_array[32445] = 32'hFFFFFFF1;
    // rom_array[32446] = 32'hFFFFFFF1;
    // rom_array[32447] = 32'hFFFFFFF1;
    // rom_array[32448] = 32'hFFFFFFF1;
    // rom_array[32449] = 32'hFFFFFFF0;
    // rom_array[32450] = 32'hFFFFFFF0;
    // rom_array[32451] = 32'hFFFFFFF0;
    // rom_array[32452] = 32'hFFFFFFF0;
    // rom_array[32453] = 32'hFFFFFFF1;
    // rom_array[32454] = 32'hFFFFFFF1;
    // rom_array[32455] = 32'hFFFFFFF1;
    // rom_array[32456] = 32'hFFFFFFF1;
    // rom_array[32457] = 32'hFFFFFFF0;
    // rom_array[32458] = 32'hFFFFFFF0;
    // rom_array[32459] = 32'hFFFFFFF0;
    // rom_array[32460] = 32'hFFFFFFF0;
    // rom_array[32461] = 32'hFFFFFFF1;
    // rom_array[32462] = 32'hFFFFFFF1;
    // rom_array[32463] = 32'hFFFFFFF1;
    // rom_array[32464] = 32'hFFFFFFF1;
    // rom_array[32465] = 32'hFFFFFFF0;
    // rom_array[32466] = 32'hFFFFFFF0;
    // rom_array[32467] = 32'hFFFFFFF0;
    // rom_array[32468] = 32'hFFFFFFF0;
    // rom_array[32469] = 32'hFFFFFFF1;
    // rom_array[32470] = 32'hFFFFFFF1;
    // rom_array[32471] = 32'hFFFFFFF1;
    // rom_array[32472] = 32'hFFFFFFF1;
    // rom_array[32473] = 32'hFFFFFFF0;
    // rom_array[32474] = 32'hFFFFFFF0;
    // rom_array[32475] = 32'hFFFFFFF0;
    // rom_array[32476] = 32'hFFFFFFF0;
    // rom_array[32477] = 32'hFFFFFFF1;
    // rom_array[32478] = 32'hFFFFFFF1;
    // rom_array[32479] = 32'hFFFFFFF1;
    // rom_array[32480] = 32'hFFFFFFF1;
    // rom_array[32481] = 32'hFFFFFFF0;
    // rom_array[32482] = 32'hFFFFFFF0;
    // rom_array[32483] = 32'hFFFFFFF0;
    // rom_array[32484] = 32'hFFFFFFF0;
    // rom_array[32485] = 32'hFFFFFFF1;
    // rom_array[32486] = 32'hFFFFFFF1;
    // rom_array[32487] = 32'hFFFFFFF1;
    // rom_array[32488] = 32'hFFFFFFF1;
    // rom_array[32489] = 32'hFFFFFFF0;
    // rom_array[32490] = 32'hFFFFFFF0;
    // rom_array[32491] = 32'hFFFFFFF0;
    // rom_array[32492] = 32'hFFFFFFF0;
    // rom_array[32493] = 32'hFFFFFFF1;
    // rom_array[32494] = 32'hFFFFFFF1;
    // rom_array[32495] = 32'hFFFFFFF1;
    // rom_array[32496] = 32'hFFFFFFF1;
    // rom_array[32497] = 32'hFFFFFFF0;
    // rom_array[32498] = 32'hFFFFFFF0;
    // rom_array[32499] = 32'hFFFFFFF0;
    // rom_array[32500] = 32'hFFFFFFF0;
    // rom_array[32501] = 32'hFFFFFFF1;
    // rom_array[32502] = 32'hFFFFFFF1;
    // rom_array[32503] = 32'hFFFFFFF1;
    // rom_array[32504] = 32'hFFFFFFF1;
    // rom_array[32505] = 32'hFFFFFFF0;
    // rom_array[32506] = 32'hFFFFFFF0;
    // rom_array[32507] = 32'hFFFFFFF0;
    // rom_array[32508] = 32'hFFFFFFF0;
    // rom_array[32509] = 32'hFFFFFFF0;
    // rom_array[32510] = 32'hFFFFFFF0;
    // rom_array[32511] = 32'hFFFFFFF1;
    // rom_array[32512] = 32'hFFFFFFF1;
    // rom_array[32513] = 32'hFFFFFFF0;
    // rom_array[32514] = 32'hFFFFFFF0;
    // rom_array[32515] = 32'hFFFFFFF0;
    // rom_array[32516] = 32'hFFFFFFF0;
    // rom_array[32517] = 32'hFFFFFFF0;
    // rom_array[32518] = 32'hFFFFFFF0;
    // rom_array[32519] = 32'hFFFFFFF1;
    // rom_array[32520] = 32'hFFFFFFF1;
    // rom_array[32521] = 32'hFFFFFFF0;
    // rom_array[32522] = 32'hFFFFFFF0;
    // rom_array[32523] = 32'hFFFFFFF0;
    // rom_array[32524] = 32'hFFFFFFF0;
    // rom_array[32525] = 32'hFFFFFFF1;
    // rom_array[32526] = 32'hFFFFFFF1;
    // rom_array[32527] = 32'hFFFFFFF1;
    // rom_array[32528] = 32'hFFFFFFF1;
    // rom_array[32529] = 32'hFFFFFFF0;
    // rom_array[32530] = 32'hFFFFFFF0;
    // rom_array[32531] = 32'hFFFFFFF0;
    // rom_array[32532] = 32'hFFFFFFF0;
    // rom_array[32533] = 32'hFFFFFFF1;
    // rom_array[32534] = 32'hFFFFFFF1;
    // rom_array[32535] = 32'hFFFFFFF1;
    // rom_array[32536] = 32'hFFFFFFF1;
    // rom_array[32537] = 32'hFFFFFFF0;
    // rom_array[32538] = 32'hFFFFFFF0;
    // rom_array[32539] = 32'hFFFFFFF0;
    // rom_array[32540] = 32'hFFFFFFF0;
    // rom_array[32541] = 32'hFFFFFFF1;
    // rom_array[32542] = 32'hFFFFFFF1;
    // rom_array[32543] = 32'hFFFFFFF1;
    // rom_array[32544] = 32'hFFFFFFF1;
    // rom_array[32545] = 32'hFFFFFFF0;
    // rom_array[32546] = 32'hFFFFFFF0;
    // rom_array[32547] = 32'hFFFFFFF0;
    // rom_array[32548] = 32'hFFFFFFF0;
    // rom_array[32549] = 32'hFFFFFFF1;
    // rom_array[32550] = 32'hFFFFFFF1;
    // rom_array[32551] = 32'hFFFFFFF1;
    // rom_array[32552] = 32'hFFFFFFF1;
    // rom_array[32553] = 32'hFFFFFFF0;
    // rom_array[32554] = 32'hFFFFFFF0;
    // rom_array[32555] = 32'hFFFFFFF0;
    // rom_array[32556] = 32'hFFFFFFF0;
    // rom_array[32557] = 32'hFFFFFFF1;
    // rom_array[32558] = 32'hFFFFFFF1;
    // rom_array[32559] = 32'hFFFFFFF1;
    // rom_array[32560] = 32'hFFFFFFF1;
    // rom_array[32561] = 32'hFFFFFFF0;
    // rom_array[32562] = 32'hFFFFFFF0;
    // rom_array[32563] = 32'hFFFFFFF0;
    // rom_array[32564] = 32'hFFFFFFF0;
    // rom_array[32565] = 32'hFFFFFFF1;
    // rom_array[32566] = 32'hFFFFFFF1;
    // rom_array[32567] = 32'hFFFFFFF1;
    // rom_array[32568] = 32'hFFFFFFF1;
    // rom_array[32569] = 32'hFFFFFFF0;
    // rom_array[32570] = 32'hFFFFFFF0;
    // rom_array[32571] = 32'hFFFFFFF1;
    // rom_array[32572] = 32'hFFFFFFF1;
    // rom_array[32573] = 32'hFFFFFFF0;
    // rom_array[32574] = 32'hFFFFFFF0;
    // rom_array[32575] = 32'hFFFFFFF1;
    // rom_array[32576] = 32'hFFFFFFF1;
    // rom_array[32577] = 32'hFFFFFFF0;
    // rom_array[32578] = 32'hFFFFFFF0;
    // rom_array[32579] = 32'hFFFFFFF1;
    // rom_array[32580] = 32'hFFFFFFF1;
    // rom_array[32581] = 32'hFFFFFFF0;
    // rom_array[32582] = 32'hFFFFFFF0;
    // rom_array[32583] = 32'hFFFFFFF1;
    // rom_array[32584] = 32'hFFFFFFF1;
    // rom_array[32585] = 32'hFFFFFFF0;
    // rom_array[32586] = 32'hFFFFFFF0;
    // rom_array[32587] = 32'hFFFFFFF1;
    // rom_array[32588] = 32'hFFFFFFF1;
    // rom_array[32589] = 32'hFFFFFFF0;
    // rom_array[32590] = 32'hFFFFFFF0;
    // rom_array[32591] = 32'hFFFFFFF1;
    // rom_array[32592] = 32'hFFFFFFF1;
    // rom_array[32593] = 32'hFFFFFFF0;
    // rom_array[32594] = 32'hFFFFFFF0;
    // rom_array[32595] = 32'hFFFFFFF1;
    // rom_array[32596] = 32'hFFFFFFF1;
    // rom_array[32597] = 32'hFFFFFFF0;
    // rom_array[32598] = 32'hFFFFFFF0;
    // rom_array[32599] = 32'hFFFFFFF1;
    // rom_array[32600] = 32'hFFFFFFF1;
    // rom_array[32601] = 32'hFFFFFFF0;
    // rom_array[32602] = 32'hFFFFFFF0;
    // rom_array[32603] = 32'hFFFFFFF0;
    // rom_array[32604] = 32'hFFFFFFF0;
    // rom_array[32605] = 32'hFFFFFFF1;
    // rom_array[32606] = 32'hFFFFFFF1;
    // rom_array[32607] = 32'hFFFFFFF1;
    // rom_array[32608] = 32'hFFFFFFF1;
    // rom_array[32609] = 32'hFFFFFFF0;
    // rom_array[32610] = 32'hFFFFFFF0;
    // rom_array[32611] = 32'hFFFFFFF0;
    // rom_array[32612] = 32'hFFFFFFF0;
    // rom_array[32613] = 32'hFFFFFFF1;
    // rom_array[32614] = 32'hFFFFFFF1;
    // rom_array[32615] = 32'hFFFFFFF1;
    // rom_array[32616] = 32'hFFFFFFF1;
    // rom_array[32617] = 32'hFFFFFFF1;
    // rom_array[32618] = 32'hFFFFFFF1;
    // rom_array[32619] = 32'hFFFFFFF1;
    // rom_array[32620] = 32'hFFFFFFF1;
    // rom_array[32621] = 32'hFFFFFFF1;
    // rom_array[32622] = 32'hFFFFFFF1;
    // rom_array[32623] = 32'hFFFFFFF1;
    // rom_array[32624] = 32'hFFFFFFF1;
    // rom_array[32625] = 32'hFFFFFFF1;
    // rom_array[32626] = 32'hFFFFFFF1;
    // rom_array[32627] = 32'hFFFFFFF1;
    // rom_array[32628] = 32'hFFFFFFF1;
    // rom_array[32629] = 32'hFFFFFFF1;
    // rom_array[32630] = 32'hFFFFFFF1;
    // rom_array[32631] = 32'hFFFFFFF1;
    // rom_array[32632] = 32'hFFFFFFF1;
    // rom_array[32633] = 32'hFFFFFFF1;
    // rom_array[32634] = 32'hFFFFFFF1;
    // rom_array[32635] = 32'hFFFFFFF1;
    // rom_array[32636] = 32'hFFFFFFF1;
    // rom_array[32637] = 32'hFFFFFFF1;
    // rom_array[32638] = 32'hFFFFFFF1;
    // rom_array[32639] = 32'hFFFFFFF1;
    // rom_array[32640] = 32'hFFFFFFF1;
    // rom_array[32641] = 32'hFFFFFFF1;
    // rom_array[32642] = 32'hFFFFFFF1;
    // rom_array[32643] = 32'hFFFFFFF1;
    // rom_array[32644] = 32'hFFFFFFF1;
    // rom_array[32645] = 32'hFFFFFFF1;
    // rom_array[32646] = 32'hFFFFFFF1;
    // rom_array[32647] = 32'hFFFFFFF1;
    // rom_array[32648] = 32'hFFFFFFF1;
    // rom_array[32649] = 32'hFFFFFFF0;
    // rom_array[32650] = 32'hFFFFFFF0;
    // rom_array[32651] = 32'hFFFFFFF1;
    // rom_array[32652] = 32'hFFFFFFF1;
    // rom_array[32653] = 32'hFFFFFFF0;
    // rom_array[32654] = 32'hFFFFFFF0;
    // rom_array[32655] = 32'hFFFFFFF1;
    // rom_array[32656] = 32'hFFFFFFF1;
    // rom_array[32657] = 32'hFFFFFFF0;
    // rom_array[32658] = 32'hFFFFFFF0;
    // rom_array[32659] = 32'hFFFFFFF1;
    // rom_array[32660] = 32'hFFFFFFF1;
    // rom_array[32661] = 32'hFFFFFFF0;
    // rom_array[32662] = 32'hFFFFFFF0;
    // rom_array[32663] = 32'hFFFFFFF1;
    // rom_array[32664] = 32'hFFFFFFF1;
    // rom_array[32665] = 32'hFFFFFFF0;
    // rom_array[32666] = 32'hFFFFFFF0;
    // rom_array[32667] = 32'hFFFFFFF0;
    // rom_array[32668] = 32'hFFFFFFF0;
    // rom_array[32669] = 32'hFFFFFFF1;
    // rom_array[32670] = 32'hFFFFFFF1;
    // rom_array[32671] = 32'hFFFFFFF1;
    // rom_array[32672] = 32'hFFFFFFF1;
    // rom_array[32673] = 32'hFFFFFFF0;
    // rom_array[32674] = 32'hFFFFFFF0;
    // rom_array[32675] = 32'hFFFFFFF0;
    // rom_array[32676] = 32'hFFFFFFF0;
    // rom_array[32677] = 32'hFFFFFFF1;
    // rom_array[32678] = 32'hFFFFFFF1;
    // rom_array[32679] = 32'hFFFFFFF1;
    // rom_array[32680] = 32'hFFFFFFF1;
    // rom_array[32681] = 32'hFFFFFFF0;
    // rom_array[32682] = 32'hFFFFFFF0;
    // rom_array[32683] = 32'hFFFFFFF1;
    // rom_array[32684] = 32'hFFFFFFF1;
    // rom_array[32685] = 32'hFFFFFFF0;
    // rom_array[32686] = 32'hFFFFFFF0;
    // rom_array[32687] = 32'hFFFFFFF1;
    // rom_array[32688] = 32'hFFFFFFF1;
    // rom_array[32689] = 32'hFFFFFFF0;
    // rom_array[32690] = 32'hFFFFFFF0;
    // rom_array[32691] = 32'hFFFFFFF1;
    // rom_array[32692] = 32'hFFFFFFF1;
    // rom_array[32693] = 32'hFFFFFFF0;
    // rom_array[32694] = 32'hFFFFFFF0;
    // rom_array[32695] = 32'hFFFFFFF1;
    // rom_array[32696] = 32'hFFFFFFF1;
    // rom_array[32697] = 32'hFFFFFFF0;
    // rom_array[32698] = 32'hFFFFFFF0;
    // rom_array[32699] = 32'hFFFFFFF0;
    // rom_array[32700] = 32'hFFFFFFF0;
    // rom_array[32701] = 32'hFFFFFFF1;
    // rom_array[32702] = 32'hFFFFFFF1;
    // rom_array[32703] = 32'hFFFFFFF1;
    // rom_array[32704] = 32'hFFFFFFF1;
    // rom_array[32705] = 32'hFFFFFFF0;
    // rom_array[32706] = 32'hFFFFFFF0;
    // rom_array[32707] = 32'hFFFFFFF0;
    // rom_array[32708] = 32'hFFFFFFF0;
    // rom_array[32709] = 32'hFFFFFFF1;
    // rom_array[32710] = 32'hFFFFFFF1;
    // rom_array[32711] = 32'hFFFFFFF1;
    // rom_array[32712] = 32'hFFFFFFF1;
    // rom_array[32713] = 32'hFFFFFFF0;
    // rom_array[32714] = 32'hFFFFFFF0;
    // rom_array[32715] = 32'hFFFFFFF0;
    // rom_array[32716] = 32'hFFFFFFF0;
    // rom_array[32717] = 32'hFFFFFFF1;
    // rom_array[32718] = 32'hFFFFFFF1;
    // rom_array[32719] = 32'hFFFFFFF1;
    // rom_array[32720] = 32'hFFFFFFF1;
    // rom_array[32721] = 32'hFFFFFFF0;
    // rom_array[32722] = 32'hFFFFFFF0;
    // rom_array[32723] = 32'hFFFFFFF0;
    // rom_array[32724] = 32'hFFFFFFF0;
    // rom_array[32725] = 32'hFFFFFFF1;
    // rom_array[32726] = 32'hFFFFFFF1;
    // rom_array[32727] = 32'hFFFFFFF1;
    // rom_array[32728] = 32'hFFFFFFF1;
    // rom_array[32729] = 32'hFFFFFFF0;
    // rom_array[32730] = 32'hFFFFFFF0;
    // rom_array[32731] = 32'hFFFFFFF1;
    // rom_array[32732] = 32'hFFFFFFF1;
    // rom_array[32733] = 32'hFFFFFFF0;
    // rom_array[32734] = 32'hFFFFFFF0;
    // rom_array[32735] = 32'hFFFFFFF1;
    // rom_array[32736] = 32'hFFFFFFF1;
    // rom_array[32737] = 32'hFFFFFFF0;
    // rom_array[32738] = 32'hFFFFFFF0;
    // rom_array[32739] = 32'hFFFFFFF1;
    // rom_array[32740] = 32'hFFFFFFF1;
    // rom_array[32741] = 32'hFFFFFFF0;
    // rom_array[32742] = 32'hFFFFFFF0;
    // rom_array[32743] = 32'hFFFFFFF1;
    // rom_array[32744] = 32'hFFFFFFF1;
    // rom_array[32745] = 32'hFFFFFFF0;
    // rom_array[32746] = 32'hFFFFFFF0;
    // rom_array[32747] = 32'hFFFFFFF1;
    // rom_array[32748] = 32'hFFFFFFF1;
    // rom_array[32749] = 32'hFFFFFFF0;
    // rom_array[32750] = 32'hFFFFFFF0;
    // rom_array[32751] = 32'hFFFFFFF1;
    // rom_array[32752] = 32'hFFFFFFF1;
    // rom_array[32753] = 32'hFFFFFFF0;
    // rom_array[32754] = 32'hFFFFFFF0;
    // rom_array[32755] = 32'hFFFFFFF1;
    // rom_array[32756] = 32'hFFFFFFF1;
    // rom_array[32757] = 32'hFFFFFFF0;
    // rom_array[32758] = 32'hFFFFFFF0;
    // rom_array[32759] = 32'hFFFFFFF1;
    // rom_array[32760] = 32'hFFFFFFF1;
    // rom_array[32761] = 32'hFFFFFFF0;
    // rom_array[32762] = 32'hFFFFFFF0;
    // rom_array[32763] = 32'hFFFFFFF1;
    // rom_array[32764] = 32'hFFFFFFF1;
    // rom_array[32765] = 32'hFFFFFFF0;
    // rom_array[32766] = 32'hFFFFFFF0;
    // rom_array[32767] = 32'hFFFFFFF1;
    // rom_array[32768] = 32'hFFFFFFF1;
    // rom_array[32769] = 32'hFFFFFFF0;
    // rom_array[32770] = 32'hFFFFFFF0;
    // rom_array[32771] = 32'hFFFFFFF1;
    // rom_array[32772] = 32'hFFFFFFF1;
    // rom_array[32773] = 32'hFFFFFFF0;
    // rom_array[32774] = 32'hFFFFFFF0;
    // rom_array[32775] = 32'hFFFFFFF1;
    // rom_array[32776] = 32'hFFFFFFF1;
    // rom_array[32777] = 32'hFFFFFFF1;
    // rom_array[32778] = 32'hFFFFFFF1;
    // rom_array[32779] = 32'hFFFFFFF1;
    // rom_array[32780] = 32'hFFFFFFF1;
    // rom_array[32781] = 32'hFFFFFFF0;
    // rom_array[32782] = 32'hFFFFFFF0;
    // rom_array[32783] = 32'hFFFFFFF0;
    // rom_array[32784] = 32'hFFFFFFF0;
    // rom_array[32785] = 32'hFFFFFFF1;
    // rom_array[32786] = 32'hFFFFFFF1;
    // rom_array[32787] = 32'hFFFFFFF1;
    // rom_array[32788] = 32'hFFFFFFF1;
    // rom_array[32789] = 32'hFFFFFFF0;
    // rom_array[32790] = 32'hFFFFFFF0;
    // rom_array[32791] = 32'hFFFFFFF0;
    // rom_array[32792] = 32'hFFFFFFF0;
    // rom_array[32793] = 32'hFFFFFFF0;
    // rom_array[32794] = 32'hFFFFFFF0;
    // rom_array[32795] = 32'hFFFFFFF1;
    // rom_array[32796] = 32'hFFFFFFF1;
    // rom_array[32797] = 32'hFFFFFFF0;
    // rom_array[32798] = 32'hFFFFFFF0;
    // rom_array[32799] = 32'hFFFFFFF1;
    // rom_array[32800] = 32'hFFFFFFF1;
    // rom_array[32801] = 32'hFFFFFFF0;
    // rom_array[32802] = 32'hFFFFFFF0;
    // rom_array[32803] = 32'hFFFFFFF1;
    // rom_array[32804] = 32'hFFFFFFF1;
    // rom_array[32805] = 32'hFFFFFFF0;
    // rom_array[32806] = 32'hFFFFFFF0;
    // rom_array[32807] = 32'hFFFFFFF1;
    // rom_array[32808] = 32'hFFFFFFF1;
    // rom_array[32809] = 32'hFFFFFFF1;
    // rom_array[32810] = 32'hFFFFFFF1;
    // rom_array[32811] = 32'hFFFFFFF1;
    // rom_array[32812] = 32'hFFFFFFF1;
    // rom_array[32813] = 32'hFFFFFFF0;
    // rom_array[32814] = 32'hFFFFFFF0;
    // rom_array[32815] = 32'hFFFFFFF0;
    // rom_array[32816] = 32'hFFFFFFF0;
    // rom_array[32817] = 32'hFFFFFFF1;
    // rom_array[32818] = 32'hFFFFFFF1;
    // rom_array[32819] = 32'hFFFFFFF1;
    // rom_array[32820] = 32'hFFFFFFF1;
    // rom_array[32821] = 32'hFFFFFFF0;
    // rom_array[32822] = 32'hFFFFFFF0;
    // rom_array[32823] = 32'hFFFFFFF0;
    // rom_array[32824] = 32'hFFFFFFF0;
    // rom_array[32825] = 32'hFFFFFFF1;
    // rom_array[32826] = 32'hFFFFFFF1;
    // rom_array[32827] = 32'hFFFFFFF1;
    // rom_array[32828] = 32'hFFFFFFF1;
    // rom_array[32829] = 32'hFFFFFFF0;
    // rom_array[32830] = 32'hFFFFFFF0;
    // rom_array[32831] = 32'hFFFFFFF0;
    // rom_array[32832] = 32'hFFFFFFF0;
    // rom_array[32833] = 32'hFFFFFFF1;
    // rom_array[32834] = 32'hFFFFFFF1;
    // rom_array[32835] = 32'hFFFFFFF1;
    // rom_array[32836] = 32'hFFFFFFF1;
    // rom_array[32837] = 32'hFFFFFFF0;
    // rom_array[32838] = 32'hFFFFFFF0;
    // rom_array[32839] = 32'hFFFFFFF0;
    // rom_array[32840] = 32'hFFFFFFF0;
    // rom_array[32841] = 32'hFFFFFFF0;
    // rom_array[32842] = 32'hFFFFFFF0;
    // rom_array[32843] = 32'hFFFFFFF1;
    // rom_array[32844] = 32'hFFFFFFF1;
    // rom_array[32845] = 32'hFFFFFFF0;
    // rom_array[32846] = 32'hFFFFFFF0;
    // rom_array[32847] = 32'hFFFFFFF1;
    // rom_array[32848] = 32'hFFFFFFF1;
    // rom_array[32849] = 32'hFFFFFFF0;
    // rom_array[32850] = 32'hFFFFFFF0;
    // rom_array[32851] = 32'hFFFFFFF1;
    // rom_array[32852] = 32'hFFFFFFF1;
    // rom_array[32853] = 32'hFFFFFFF0;
    // rom_array[32854] = 32'hFFFFFFF0;
    // rom_array[32855] = 32'hFFFFFFF1;
    // rom_array[32856] = 32'hFFFFFFF1;
    // rom_array[32857] = 32'hFFFFFFF0;
    // rom_array[32858] = 32'hFFFFFFF0;
    // rom_array[32859] = 32'hFFFFFFF1;
    // rom_array[32860] = 32'hFFFFFFF1;
    // rom_array[32861] = 32'hFFFFFFF0;
    // rom_array[32862] = 32'hFFFFFFF0;
    // rom_array[32863] = 32'hFFFFFFF1;
    // rom_array[32864] = 32'hFFFFFFF1;
    // rom_array[32865] = 32'hFFFFFFF0;
    // rom_array[32866] = 32'hFFFFFFF0;
    // rom_array[32867] = 32'hFFFFFFF1;
    // rom_array[32868] = 32'hFFFFFFF1;
    // rom_array[32869] = 32'hFFFFFFF0;
    // rom_array[32870] = 32'hFFFFFFF0;
    // rom_array[32871] = 32'hFFFFFFF1;
    // rom_array[32872] = 32'hFFFFFFF1;
    // rom_array[32873] = 32'hFFFFFFF0;
    // rom_array[32874] = 32'hFFFFFFF0;
    // rom_array[32875] = 32'hFFFFFFF1;
    // rom_array[32876] = 32'hFFFFFFF1;
    // rom_array[32877] = 32'hFFFFFFF1;
    // rom_array[32878] = 32'hFFFFFFF1;
    // rom_array[32879] = 32'hFFFFFFF1;
    // rom_array[32880] = 32'hFFFFFFF1;
    // rom_array[32881] = 32'hFFFFFFF0;
    // rom_array[32882] = 32'hFFFFFFF0;
    // rom_array[32883] = 32'hFFFFFFF1;
    // rom_array[32884] = 32'hFFFFFFF1;
    // rom_array[32885] = 32'hFFFFFFF1;
    // rom_array[32886] = 32'hFFFFFFF1;
    // rom_array[32887] = 32'hFFFFFFF1;
    // rom_array[32888] = 32'hFFFFFFF1;
    // rom_array[32889] = 32'hFFFFFFF0;
    // rom_array[32890] = 32'hFFFFFFF0;
    // rom_array[32891] = 32'hFFFFFFF0;
    // rom_array[32892] = 32'hFFFFFFF0;
    // rom_array[32893] = 32'hFFFFFFF1;
    // rom_array[32894] = 32'hFFFFFFF1;
    // rom_array[32895] = 32'hFFFFFFF1;
    // rom_array[32896] = 32'hFFFFFFF1;
    // rom_array[32897] = 32'hFFFFFFF0;
    // rom_array[32898] = 32'hFFFFFFF0;
    // rom_array[32899] = 32'hFFFFFFF0;
    // rom_array[32900] = 32'hFFFFFFF0;
    // rom_array[32901] = 32'hFFFFFFF1;
    // rom_array[32902] = 32'hFFFFFFF1;
    // rom_array[32903] = 32'hFFFFFFF1;
    // rom_array[32904] = 32'hFFFFFFF1;
    // rom_array[32905] = 32'hFFFFFFF0;
    // rom_array[32906] = 32'hFFFFFFF0;
    // rom_array[32907] = 32'hFFFFFFF1;
    // rom_array[32908] = 32'hFFFFFFF1;
    // rom_array[32909] = 32'hFFFFFFF0;
    // rom_array[32910] = 32'hFFFFFFF0;
    // rom_array[32911] = 32'hFFFFFFF1;
    // rom_array[32912] = 32'hFFFFFFF1;
    // rom_array[32913] = 32'hFFFFFFF0;
    // rom_array[32914] = 32'hFFFFFFF0;
    // rom_array[32915] = 32'hFFFFFFF1;
    // rom_array[32916] = 32'hFFFFFFF1;
    // rom_array[32917] = 32'hFFFFFFF0;
    // rom_array[32918] = 32'hFFFFFFF0;
    // rom_array[32919] = 32'hFFFFFFF1;
    // rom_array[32920] = 32'hFFFFFFF1;
    // rom_array[32921] = 32'hFFFFFFF0;
    // rom_array[32922] = 32'hFFFFFFF0;
    // rom_array[32923] = 32'hFFFFFFF0;
    // rom_array[32924] = 32'hFFFFFFF0;
    // rom_array[32925] = 32'hFFFFFFF1;
    // rom_array[32926] = 32'hFFFFFFF1;
    // rom_array[32927] = 32'hFFFFFFF1;
    // rom_array[32928] = 32'hFFFFFFF1;
    // rom_array[32929] = 32'hFFFFFFF0;
    // rom_array[32930] = 32'hFFFFFFF0;
    // rom_array[32931] = 32'hFFFFFFF0;
    // rom_array[32932] = 32'hFFFFFFF0;
    // rom_array[32933] = 32'hFFFFFFF1;
    // rom_array[32934] = 32'hFFFFFFF1;
    // rom_array[32935] = 32'hFFFFFFF1;
    // rom_array[32936] = 32'hFFFFFFF1;
    // rom_array[32937] = 32'hFFFFFFF0;
    // rom_array[32938] = 32'hFFFFFFF0;
    // rom_array[32939] = 32'hFFFFFFF0;
    // rom_array[32940] = 32'hFFFFFFF0;
    // rom_array[32941] = 32'hFFFFFFF1;
    // rom_array[32942] = 32'hFFFFFFF1;
    // rom_array[32943] = 32'hFFFFFFF1;
    // rom_array[32944] = 32'hFFFFFFF1;
    // rom_array[32945] = 32'hFFFFFFF0;
    // rom_array[32946] = 32'hFFFFFFF0;
    // rom_array[32947] = 32'hFFFFFFF0;
    // rom_array[32948] = 32'hFFFFFFF0;
    // rom_array[32949] = 32'hFFFFFFF1;
    // rom_array[32950] = 32'hFFFFFFF1;
    // rom_array[32951] = 32'hFFFFFFF1;
    // rom_array[32952] = 32'hFFFFFFF1;
    // rom_array[32953] = 32'hFFFFFFF0;
    // rom_array[32954] = 32'hFFFFFFF0;
    // rom_array[32955] = 32'hFFFFFFF1;
    // rom_array[32956] = 32'hFFFFFFF1;
    // rom_array[32957] = 32'hFFFFFFF0;
    // rom_array[32958] = 32'hFFFFFFF0;
    // rom_array[32959] = 32'hFFFFFFF1;
    // rom_array[32960] = 32'hFFFFFFF1;
    // rom_array[32961] = 32'hFFFFFFF0;
    // rom_array[32962] = 32'hFFFFFFF0;
    // rom_array[32963] = 32'hFFFFFFF1;
    // rom_array[32964] = 32'hFFFFFFF1;
    // rom_array[32965] = 32'hFFFFFFF0;
    // rom_array[32966] = 32'hFFFFFFF0;
    // rom_array[32967] = 32'hFFFFFFF1;
    // rom_array[32968] = 32'hFFFFFFF1;
    // rom_array[32969] = 32'hFFFFFFF0;
    // rom_array[32970] = 32'hFFFFFFF0;
    // rom_array[32971] = 32'hFFFFFFF1;
    // rom_array[32972] = 32'hFFFFFFF1;
    // rom_array[32973] = 32'hFFFFFFF0;
    // rom_array[32974] = 32'hFFFFFFF0;
    // rom_array[32975] = 32'hFFFFFFF1;
    // rom_array[32976] = 32'hFFFFFFF1;
    // rom_array[32977] = 32'hFFFFFFF0;
    // rom_array[32978] = 32'hFFFFFFF0;
    // rom_array[32979] = 32'hFFFFFFF1;
    // rom_array[32980] = 32'hFFFFFFF1;
    // rom_array[32981] = 32'hFFFFFFF0;
    // rom_array[32982] = 32'hFFFFFFF0;
    // rom_array[32983] = 32'hFFFFFFF1;
    // rom_array[32984] = 32'hFFFFFFF1;
    // rom_array[32985] = 32'hFFFFFFF1;
    // rom_array[32986] = 32'hFFFFFFF1;
    // rom_array[32987] = 32'hFFFFFFF1;
    // rom_array[32988] = 32'hFFFFFFF1;
    // rom_array[32989] = 32'hFFFFFFF1;
    // rom_array[32990] = 32'hFFFFFFF1;
    // rom_array[32991] = 32'hFFFFFFF1;
    // rom_array[32992] = 32'hFFFFFFF1;
    // rom_array[32993] = 32'hFFFFFFF1;
    // rom_array[32994] = 32'hFFFFFFF1;
    // rom_array[32995] = 32'hFFFFFFF1;
    // rom_array[32996] = 32'hFFFFFFF1;
    // rom_array[32997] = 32'hFFFFFFF1;
    // rom_array[32998] = 32'hFFFFFFF1;
    // rom_array[32999] = 32'hFFFFFFF1;
    // rom_array[33000] = 32'hFFFFFFF1;
    // rom_array[33001] = 32'hFFFFFFF0;
    // rom_array[33002] = 32'hFFFFFFF0;
    // rom_array[33003] = 32'hFFFFFFF0;
    // rom_array[33004] = 32'hFFFFFFF0;
    // rom_array[33005] = 32'hFFFFFFF1;
    // rom_array[33006] = 32'hFFFFFFF1;
    // rom_array[33007] = 32'hFFFFFFF1;
    // rom_array[33008] = 32'hFFFFFFF1;
    // rom_array[33009] = 32'hFFFFFFF0;
    // rom_array[33010] = 32'hFFFFFFF0;
    // rom_array[33011] = 32'hFFFFFFF0;
    // rom_array[33012] = 32'hFFFFFFF0;
    // rom_array[33013] = 32'hFFFFFFF1;
    // rom_array[33014] = 32'hFFFFFFF1;
    // rom_array[33015] = 32'hFFFFFFF1;
    // rom_array[33016] = 32'hFFFFFFF1;
    // rom_array[33017] = 32'hFFFFFFF1;
    // rom_array[33018] = 32'hFFFFFFF1;
    // rom_array[33019] = 32'hFFFFFFF1;
    // rom_array[33020] = 32'hFFFFFFF1;
    // rom_array[33021] = 32'hFFFFFFF1;
    // rom_array[33022] = 32'hFFFFFFF1;
    // rom_array[33023] = 32'hFFFFFFF1;
    // rom_array[33024] = 32'hFFFFFFF1;
    // rom_array[33025] = 32'hFFFFFFF1;
    // rom_array[33026] = 32'hFFFFFFF1;
    // rom_array[33027] = 32'hFFFFFFF1;
    // rom_array[33028] = 32'hFFFFFFF1;
    // rom_array[33029] = 32'hFFFFFFF1;
    // rom_array[33030] = 32'hFFFFFFF1;
    // rom_array[33031] = 32'hFFFFFFF1;
    // rom_array[33032] = 32'hFFFFFFF1;
    // rom_array[33033] = 32'hFFFFFFF0;
    // rom_array[33034] = 32'hFFFFFFF0;
    // rom_array[33035] = 32'hFFFFFFF0;
    // rom_array[33036] = 32'hFFFFFFF0;
    // rom_array[33037] = 32'hFFFFFFF1;
    // rom_array[33038] = 32'hFFFFFFF1;
    // rom_array[33039] = 32'hFFFFFFF1;
    // rom_array[33040] = 32'hFFFFFFF1;
    // rom_array[33041] = 32'hFFFFFFF0;
    // rom_array[33042] = 32'hFFFFFFF0;
    // rom_array[33043] = 32'hFFFFFFF0;
    // rom_array[33044] = 32'hFFFFFFF0;
    // rom_array[33045] = 32'hFFFFFFF1;
    // rom_array[33046] = 32'hFFFFFFF1;
    // rom_array[33047] = 32'hFFFFFFF1;
    // rom_array[33048] = 32'hFFFFFFF1;
    // rom_array[33049] = 32'hFFFFFFF0;
    // rom_array[33050] = 32'hFFFFFFF0;
    // rom_array[33051] = 32'hFFFFFFF0;
    // rom_array[33052] = 32'hFFFFFFF0;
    // rom_array[33053] = 32'hFFFFFFF1;
    // rom_array[33054] = 32'hFFFFFFF1;
    // rom_array[33055] = 32'hFFFFFFF1;
    // rom_array[33056] = 32'hFFFFFFF1;
    // rom_array[33057] = 32'hFFFFFFF0;
    // rom_array[33058] = 32'hFFFFFFF0;
    // rom_array[33059] = 32'hFFFFFFF0;
    // rom_array[33060] = 32'hFFFFFFF0;
    // rom_array[33061] = 32'hFFFFFFF1;
    // rom_array[33062] = 32'hFFFFFFF1;
    // rom_array[33063] = 32'hFFFFFFF1;
    // rom_array[33064] = 32'hFFFFFFF1;
    // rom_array[33065] = 32'hFFFFFFF1;
    // rom_array[33066] = 32'hFFFFFFF1;
    // rom_array[33067] = 32'hFFFFFFF1;
    // rom_array[33068] = 32'hFFFFFFF1;
    // rom_array[33069] = 32'hFFFFFFF1;
    // rom_array[33070] = 32'hFFFFFFF1;
    // rom_array[33071] = 32'hFFFFFFF1;
    // rom_array[33072] = 32'hFFFFFFF1;
    // rom_array[33073] = 32'hFFFFFFF1;
    // rom_array[33074] = 32'hFFFFFFF1;
    // rom_array[33075] = 32'hFFFFFFF1;
    // rom_array[33076] = 32'hFFFFFFF1;
    // rom_array[33077] = 32'hFFFFFFF1;
    // rom_array[33078] = 32'hFFFFFFF1;
    // rom_array[33079] = 32'hFFFFFFF1;
    // rom_array[33080] = 32'hFFFFFFF1;
    // rom_array[33081] = 32'hFFFFFFF1;
    // rom_array[33082] = 32'hFFFFFFF1;
    // rom_array[33083] = 32'hFFFFFFF1;
    // rom_array[33084] = 32'hFFFFFFF1;
    // rom_array[33085] = 32'hFFFFFFF1;
    // rom_array[33086] = 32'hFFFFFFF1;
    // rom_array[33087] = 32'hFFFFFFF1;
    // rom_array[33088] = 32'hFFFFFFF1;
    // rom_array[33089] = 32'hFFFFFFF1;
    // rom_array[33090] = 32'hFFFFFFF1;
    // rom_array[33091] = 32'hFFFFFFF1;
    // rom_array[33092] = 32'hFFFFFFF1;
    // rom_array[33093] = 32'hFFFFFFF1;
    // rom_array[33094] = 32'hFFFFFFF1;
    // rom_array[33095] = 32'hFFFFFFF1;
    // rom_array[33096] = 32'hFFFFFFF1;
    // rom_array[33097] = 32'hFFFFFFF1;
    // rom_array[33098] = 32'hFFFFFFF1;
    // rom_array[33099] = 32'hFFFFFFF1;
    // rom_array[33100] = 32'hFFFFFFF1;
    // rom_array[33101] = 32'hFFFFFFF0;
    // rom_array[33102] = 32'hFFFFFFF0;
    // rom_array[33103] = 32'hFFFFFFF1;
    // rom_array[33104] = 32'hFFFFFFF1;
    // rom_array[33105] = 32'hFFFFFFF1;
    // rom_array[33106] = 32'hFFFFFFF1;
    // rom_array[33107] = 32'hFFFFFFF1;
    // rom_array[33108] = 32'hFFFFFFF1;
    // rom_array[33109] = 32'hFFFFFFF0;
    // rom_array[33110] = 32'hFFFFFFF0;
    // rom_array[33111] = 32'hFFFFFFF1;
    // rom_array[33112] = 32'hFFFFFFF1;
    // rom_array[33113] = 32'hFFFFFFF1;
    // rom_array[33114] = 32'hFFFFFFF1;
    // rom_array[33115] = 32'hFFFFFFF1;
    // rom_array[33116] = 32'hFFFFFFF1;
    // rom_array[33117] = 32'hFFFFFFF0;
    // rom_array[33118] = 32'hFFFFFFF0;
    // rom_array[33119] = 32'hFFFFFFF0;
    // rom_array[33120] = 32'hFFFFFFF0;
    // rom_array[33121] = 32'hFFFFFFF1;
    // rom_array[33122] = 32'hFFFFFFF1;
    // rom_array[33123] = 32'hFFFFFFF1;
    // rom_array[33124] = 32'hFFFFFFF1;
    // rom_array[33125] = 32'hFFFFFFF0;
    // rom_array[33126] = 32'hFFFFFFF0;
    // rom_array[33127] = 32'hFFFFFFF0;
    // rom_array[33128] = 32'hFFFFFFF0;
    // rom_array[33129] = 32'hFFFFFFF0;
    // rom_array[33130] = 32'hFFFFFFF0;
    // rom_array[33131] = 32'hFFFFFFF1;
    // rom_array[33132] = 32'hFFFFFFF1;
    // rom_array[33133] = 32'hFFFFFFF0;
    // rom_array[33134] = 32'hFFFFFFF0;
    // rom_array[33135] = 32'hFFFFFFF1;
    // rom_array[33136] = 32'hFFFFFFF1;
    // rom_array[33137] = 32'hFFFFFFF0;
    // rom_array[33138] = 32'hFFFFFFF0;
    // rom_array[33139] = 32'hFFFFFFF1;
    // rom_array[33140] = 32'hFFFFFFF1;
    // rom_array[33141] = 32'hFFFFFFF0;
    // rom_array[33142] = 32'hFFFFFFF0;
    // rom_array[33143] = 32'hFFFFFFF1;
    // rom_array[33144] = 32'hFFFFFFF1;
    // rom_array[33145] = 32'hFFFFFFF1;
    // rom_array[33146] = 32'hFFFFFFF1;
    // rom_array[33147] = 32'hFFFFFFF1;
    // rom_array[33148] = 32'hFFFFFFF1;
    // rom_array[33149] = 32'hFFFFFFF0;
    // rom_array[33150] = 32'hFFFFFFF0;
    // rom_array[33151] = 32'hFFFFFFF0;
    // rom_array[33152] = 32'hFFFFFFF0;
    // rom_array[33153] = 32'hFFFFFFF1;
    // rom_array[33154] = 32'hFFFFFFF1;
    // rom_array[33155] = 32'hFFFFFFF1;
    // rom_array[33156] = 32'hFFFFFFF1;
    // rom_array[33157] = 32'hFFFFFFF0;
    // rom_array[33158] = 32'hFFFFFFF0;
    // rom_array[33159] = 32'hFFFFFFF0;
    // rom_array[33160] = 32'hFFFFFFF0;
    // rom_array[33161] = 32'hFFFFFFF1;
    // rom_array[33162] = 32'hFFFFFFF1;
    // rom_array[33163] = 32'hFFFFFFF1;
    // rom_array[33164] = 32'hFFFFFFF1;
    // rom_array[33165] = 32'hFFFFFFF0;
    // rom_array[33166] = 32'hFFFFFFF0;
    // rom_array[33167] = 32'hFFFFFFF0;
    // rom_array[33168] = 32'hFFFFFFF0;
    // rom_array[33169] = 32'hFFFFFFF1;
    // rom_array[33170] = 32'hFFFFFFF1;
    // rom_array[33171] = 32'hFFFFFFF1;
    // rom_array[33172] = 32'hFFFFFFF1;
    // rom_array[33173] = 32'hFFFFFFF0;
    // rom_array[33174] = 32'hFFFFFFF0;
    // rom_array[33175] = 32'hFFFFFFF0;
    // rom_array[33176] = 32'hFFFFFFF0;
    // rom_array[33177] = 32'hFFFFFFF0;
    // rom_array[33178] = 32'hFFFFFFF0;
    // rom_array[33179] = 32'hFFFFFFF1;
    // rom_array[33180] = 32'hFFFFFFF1;
    // rom_array[33181] = 32'hFFFFFFF0;
    // rom_array[33182] = 32'hFFFFFFF0;
    // rom_array[33183] = 32'hFFFFFFF1;
    // rom_array[33184] = 32'hFFFFFFF1;
    // rom_array[33185] = 32'hFFFFFFF0;
    // rom_array[33186] = 32'hFFFFFFF0;
    // rom_array[33187] = 32'hFFFFFFF1;
    // rom_array[33188] = 32'hFFFFFFF1;
    // rom_array[33189] = 32'hFFFFFFF0;
    // rom_array[33190] = 32'hFFFFFFF0;
    // rom_array[33191] = 32'hFFFFFFF1;
    // rom_array[33192] = 32'hFFFFFFF1;
    // rom_array[33193] = 32'hFFFFFFF0;
    // rom_array[33194] = 32'hFFFFFFF0;
    // rom_array[33195] = 32'hFFFFFFF1;
    // rom_array[33196] = 32'hFFFFFFF1;
    // rom_array[33197] = 32'hFFFFFFF0;
    // rom_array[33198] = 32'hFFFFFFF0;
    // rom_array[33199] = 32'hFFFFFFF0;
    // rom_array[33200] = 32'hFFFFFFF0;
    // rom_array[33201] = 32'hFFFFFFF0;
    // rom_array[33202] = 32'hFFFFFFF0;
    // rom_array[33203] = 32'hFFFFFFF1;
    // rom_array[33204] = 32'hFFFFFFF1;
    // rom_array[33205] = 32'hFFFFFFF0;
    // rom_array[33206] = 32'hFFFFFFF0;
    // rom_array[33207] = 32'hFFFFFFF0;
    // rom_array[33208] = 32'hFFFFFFF0;
    // rom_array[33209] = 32'hFFFFFFF1;
    // rom_array[33210] = 32'hFFFFFFF1;
    // rom_array[33211] = 32'hFFFFFFF1;
    // rom_array[33212] = 32'hFFFFFFF1;
    // rom_array[33213] = 32'hFFFFFFF0;
    // rom_array[33214] = 32'hFFFFFFF0;
    // rom_array[33215] = 32'hFFFFFFF0;
    // rom_array[33216] = 32'hFFFFFFF0;
    // rom_array[33217] = 32'hFFFFFFF1;
    // rom_array[33218] = 32'hFFFFFFF1;
    // rom_array[33219] = 32'hFFFFFFF1;
    // rom_array[33220] = 32'hFFFFFFF1;
    // rom_array[33221] = 32'hFFFFFFF0;
    // rom_array[33222] = 32'hFFFFFFF0;
    // rom_array[33223] = 32'hFFFFFFF0;
    // rom_array[33224] = 32'hFFFFFFF0;
    // rom_array[33225] = 32'hFFFFFFF1;
    // rom_array[33226] = 32'hFFFFFFF1;
    // rom_array[33227] = 32'hFFFFFFF1;
    // rom_array[33228] = 32'hFFFFFFF1;
    // rom_array[33229] = 32'hFFFFFFF0;
    // rom_array[33230] = 32'hFFFFFFF0;
    // rom_array[33231] = 32'hFFFFFFF0;
    // rom_array[33232] = 32'hFFFFFFF0;
    // rom_array[33233] = 32'hFFFFFFF1;
    // rom_array[33234] = 32'hFFFFFFF1;
    // rom_array[33235] = 32'hFFFFFFF1;
    // rom_array[33236] = 32'hFFFFFFF1;
    // rom_array[33237] = 32'hFFFFFFF0;
    // rom_array[33238] = 32'hFFFFFFF0;
    // rom_array[33239] = 32'hFFFFFFF0;
    // rom_array[33240] = 32'hFFFFFFF0;
    // rom_array[33241] = 32'hFFFFFFF1;
    // rom_array[33242] = 32'hFFFFFFF1;
    // rom_array[33243] = 32'hFFFFFFF1;
    // rom_array[33244] = 32'hFFFFFFF1;
    // rom_array[33245] = 32'hFFFFFFF0;
    // rom_array[33246] = 32'hFFFFFFF0;
    // rom_array[33247] = 32'hFFFFFFF0;
    // rom_array[33248] = 32'hFFFFFFF0;
    // rom_array[33249] = 32'hFFFFFFF1;
    // rom_array[33250] = 32'hFFFFFFF1;
    // rom_array[33251] = 32'hFFFFFFF1;
    // rom_array[33252] = 32'hFFFFFFF1;
    // rom_array[33253] = 32'hFFFFFFF0;
    // rom_array[33254] = 32'hFFFFFFF0;
    // rom_array[33255] = 32'hFFFFFFF0;
    // rom_array[33256] = 32'hFFFFFFF0;
    // rom_array[33257] = 32'hFFFFFFF1;
    // rom_array[33258] = 32'hFFFFFFF1;
    // rom_array[33259] = 32'hFFFFFFF1;
    // rom_array[33260] = 32'hFFFFFFF1;
    // rom_array[33261] = 32'hFFFFFFF1;
    // rom_array[33262] = 32'hFFFFFFF1;
    // rom_array[33263] = 32'hFFFFFFF1;
    // rom_array[33264] = 32'hFFFFFFF1;
    // rom_array[33265] = 32'hFFFFFFF1;
    // rom_array[33266] = 32'hFFFFFFF1;
    // rom_array[33267] = 32'hFFFFFFF1;
    // rom_array[33268] = 32'hFFFFFFF1;
    // rom_array[33269] = 32'hFFFFFFF1;
    // rom_array[33270] = 32'hFFFFFFF1;
    // rom_array[33271] = 32'hFFFFFFF1;
    // rom_array[33272] = 32'hFFFFFFF1;
    // rom_array[33273] = 32'hFFFFFFF1;
    // rom_array[33274] = 32'hFFFFFFF1;
    // rom_array[33275] = 32'hFFFFFFF1;
    // rom_array[33276] = 32'hFFFFFFF1;
    // rom_array[33277] = 32'hFFFFFFF0;
    // rom_array[33278] = 32'hFFFFFFF0;
    // rom_array[33279] = 32'hFFFFFFF0;
    // rom_array[33280] = 32'hFFFFFFF0;
    // rom_array[33281] = 32'hFFFFFFF1;
    // rom_array[33282] = 32'hFFFFFFF1;
    // rom_array[33283] = 32'hFFFFFFF1;
    // rom_array[33284] = 32'hFFFFFFF1;
    // rom_array[33285] = 32'hFFFFFFF0;
    // rom_array[33286] = 32'hFFFFFFF0;
    // rom_array[33287] = 32'hFFFFFFF0;
    // rom_array[33288] = 32'hFFFFFFF0;
    // rom_array[33289] = 32'hFFFFFFF1;
    // rom_array[33290] = 32'hFFFFFFF1;
    // rom_array[33291] = 32'hFFFFFFF1;
    // rom_array[33292] = 32'hFFFFFFF1;
    // rom_array[33293] = 32'hFFFFFFF1;
    // rom_array[33294] = 32'hFFFFFFF1;
    // rom_array[33295] = 32'hFFFFFFF1;
    // rom_array[33296] = 32'hFFFFFFF1;
    // rom_array[33297] = 32'hFFFFFFF1;
    // rom_array[33298] = 32'hFFFFFFF1;
    // rom_array[33299] = 32'hFFFFFFF1;
    // rom_array[33300] = 32'hFFFFFFF1;
    // rom_array[33301] = 32'hFFFFFFF1;
    // rom_array[33302] = 32'hFFFFFFF1;
    // rom_array[33303] = 32'hFFFFFFF1;
    // rom_array[33304] = 32'hFFFFFFF1;
    // rom_array[33305] = 32'hFFFFFFF1;
    // rom_array[33306] = 32'hFFFFFFF1;
    // rom_array[33307] = 32'hFFFFFFF1;
    // rom_array[33308] = 32'hFFFFFFF1;
    // rom_array[33309] = 32'hFFFFFFF0;
    // rom_array[33310] = 32'hFFFFFFF0;
    // rom_array[33311] = 32'hFFFFFFF0;
    // rom_array[33312] = 32'hFFFFFFF0;
    // rom_array[33313] = 32'hFFFFFFF1;
    // rom_array[33314] = 32'hFFFFFFF1;
    // rom_array[33315] = 32'hFFFFFFF1;
    // rom_array[33316] = 32'hFFFFFFF1;
    // rom_array[33317] = 32'hFFFFFFF0;
    // rom_array[33318] = 32'hFFFFFFF0;
    // rom_array[33319] = 32'hFFFFFFF0;
    // rom_array[33320] = 32'hFFFFFFF0;
    // rom_array[33321] = 32'hFFFFFFF1;
    // rom_array[33322] = 32'hFFFFFFF1;
    // rom_array[33323] = 32'hFFFFFFF1;
    // rom_array[33324] = 32'hFFFFFFF1;
    // rom_array[33325] = 32'hFFFFFFF0;
    // rom_array[33326] = 32'hFFFFFFF0;
    // rom_array[33327] = 32'hFFFFFFF0;
    // rom_array[33328] = 32'hFFFFFFF0;
    // rom_array[33329] = 32'hFFFFFFF1;
    // rom_array[33330] = 32'hFFFFFFF1;
    // rom_array[33331] = 32'hFFFFFFF1;
    // rom_array[33332] = 32'hFFFFFFF1;
    // rom_array[33333] = 32'hFFFFFFF0;
    // rom_array[33334] = 32'hFFFFFFF0;
    // rom_array[33335] = 32'hFFFFFFF0;
    // rom_array[33336] = 32'hFFFFFFF0;
    // rom_array[33337] = 32'hFFFFFFF1;
    // rom_array[33338] = 32'hFFFFFFF1;
    // rom_array[33339] = 32'hFFFFFFF1;
    // rom_array[33340] = 32'hFFFFFFF1;
    // rom_array[33341] = 32'hFFFFFFF1;
    // rom_array[33342] = 32'hFFFFFFF1;
    // rom_array[33343] = 32'hFFFFFFF1;
    // rom_array[33344] = 32'hFFFFFFF1;
    // rom_array[33345] = 32'hFFFFFFF1;
    // rom_array[33346] = 32'hFFFFFFF1;
    // rom_array[33347] = 32'hFFFFFFF1;
    // rom_array[33348] = 32'hFFFFFFF1;
    // rom_array[33349] = 32'hFFFFFFF1;
    // rom_array[33350] = 32'hFFFFFFF1;
    // rom_array[33351] = 32'hFFFFFFF1;
    // rom_array[33352] = 32'hFFFFFFF1;
    // rom_array[33353] = 32'hFFFFFFF1;
    // rom_array[33354] = 32'hFFFFFFF1;
    // rom_array[33355] = 32'hFFFFFFF1;
    // rom_array[33356] = 32'hFFFFFFF1;
    // rom_array[33357] = 32'hFFFFFFF0;
    // rom_array[33358] = 32'hFFFFFFF0;
    // rom_array[33359] = 32'hFFFFFFF0;
    // rom_array[33360] = 32'hFFFFFFF0;
    // rom_array[33361] = 32'hFFFFFFF1;
    // rom_array[33362] = 32'hFFFFFFF1;
    // rom_array[33363] = 32'hFFFFFFF1;
    // rom_array[33364] = 32'hFFFFFFF1;
    // rom_array[33365] = 32'hFFFFFFF0;
    // rom_array[33366] = 32'hFFFFFFF0;
    // rom_array[33367] = 32'hFFFFFFF0;
    // rom_array[33368] = 32'hFFFFFFF0;
    // rom_array[33369] = 32'hFFFFFFF0;
    // rom_array[33370] = 32'hFFFFFFF0;
    // rom_array[33371] = 32'hFFFFFFF1;
    // rom_array[33372] = 32'hFFFFFFF1;
    // rom_array[33373] = 32'hFFFFFFF0;
    // rom_array[33374] = 32'hFFFFFFF0;
    // rom_array[33375] = 32'hFFFFFFF1;
    // rom_array[33376] = 32'hFFFFFFF1;
    // rom_array[33377] = 32'hFFFFFFF0;
    // rom_array[33378] = 32'hFFFFFFF0;
    // rom_array[33379] = 32'hFFFFFFF1;
    // rom_array[33380] = 32'hFFFFFFF1;
    // rom_array[33381] = 32'hFFFFFFF0;
    // rom_array[33382] = 32'hFFFFFFF0;
    // rom_array[33383] = 32'hFFFFFFF1;
    // rom_array[33384] = 32'hFFFFFFF1;
    // rom_array[33385] = 32'hFFFFFFF1;
    // rom_array[33386] = 32'hFFFFFFF1;
    // rom_array[33387] = 32'hFFFFFFF1;
    // rom_array[33388] = 32'hFFFFFFF1;
    // rom_array[33389] = 32'hFFFFFFF1;
    // rom_array[33390] = 32'hFFFFFFF1;
    // rom_array[33391] = 32'hFFFFFFF1;
    // rom_array[33392] = 32'hFFFFFFF1;
    // rom_array[33393] = 32'hFFFFFFF1;
    // rom_array[33394] = 32'hFFFFFFF1;
    // rom_array[33395] = 32'hFFFFFFF1;
    // rom_array[33396] = 32'hFFFFFFF1;
    // rom_array[33397] = 32'hFFFFFFF1;
    // rom_array[33398] = 32'hFFFFFFF1;
    // rom_array[33399] = 32'hFFFFFFF1;
    // rom_array[33400] = 32'hFFFFFFF1;
    // rom_array[33401] = 32'hFFFFFFF0;
    // rom_array[33402] = 32'hFFFFFFF0;
    // rom_array[33403] = 32'hFFFFFFF1;
    // rom_array[33404] = 32'hFFFFFFF1;
    // rom_array[33405] = 32'hFFFFFFF0;
    // rom_array[33406] = 32'hFFFFFFF0;
    // rom_array[33407] = 32'hFFFFFFF1;
    // rom_array[33408] = 32'hFFFFFFF1;
    // rom_array[33409] = 32'hFFFFFFF0;
    // rom_array[33410] = 32'hFFFFFFF0;
    // rom_array[33411] = 32'hFFFFFFF1;
    // rom_array[33412] = 32'hFFFFFFF1;
    // rom_array[33413] = 32'hFFFFFFF0;
    // rom_array[33414] = 32'hFFFFFFF0;
    // rom_array[33415] = 32'hFFFFFFF1;
    // rom_array[33416] = 32'hFFFFFFF1;
    // rom_array[33417] = 32'hFFFFFFF1;
    // rom_array[33418] = 32'hFFFFFFF1;
    // rom_array[33419] = 32'hFFFFFFF1;
    // rom_array[33420] = 32'hFFFFFFF1;
    // rom_array[33421] = 32'hFFFFFFF1;
    // rom_array[33422] = 32'hFFFFFFF1;
    // rom_array[33423] = 32'hFFFFFFF1;
    // rom_array[33424] = 32'hFFFFFFF1;
    // rom_array[33425] = 32'hFFFFFFF1;
    // rom_array[33426] = 32'hFFFFFFF1;
    // rom_array[33427] = 32'hFFFFFFF1;
    // rom_array[33428] = 32'hFFFFFFF1;
    // rom_array[33429] = 32'hFFFFFFF1;
    // rom_array[33430] = 32'hFFFFFFF1;
    // rom_array[33431] = 32'hFFFFFFF1;
    // rom_array[33432] = 32'hFFFFFFF1;
    // rom_array[33433] = 32'hFFFFFFF1;
    // rom_array[33434] = 32'hFFFFFFF1;
    // rom_array[33435] = 32'hFFFFFFF1;
    // rom_array[33436] = 32'hFFFFFFF1;
    // rom_array[33437] = 32'hFFFFFFF1;
    // rom_array[33438] = 32'hFFFFFFF1;
    // rom_array[33439] = 32'hFFFFFFF1;
    // rom_array[33440] = 32'hFFFFFFF1;
    // rom_array[33441] = 32'hFFFFFFF1;
    // rom_array[33442] = 32'hFFFFFFF1;
    // rom_array[33443] = 32'hFFFFFFF1;
    // rom_array[33444] = 32'hFFFFFFF1;
    // rom_array[33445] = 32'hFFFFFFF1;
    // rom_array[33446] = 32'hFFFFFFF1;
    // rom_array[33447] = 32'hFFFFFFF1;
    // rom_array[33448] = 32'hFFFFFFF1;
    // rom_array[33449] = 32'hFFFFFFF1;
    // rom_array[33450] = 32'hFFFFFFF1;
    // rom_array[33451] = 32'hFFFFFFF1;
    // rom_array[33452] = 32'hFFFFFFF1;
    // rom_array[33453] = 32'hFFFFFFF1;
    // rom_array[33454] = 32'hFFFFFFF1;
    // rom_array[33455] = 32'hFFFFFFF1;
    // rom_array[33456] = 32'hFFFFFFF1;
    // rom_array[33457] = 32'hFFFFFFF1;
    // rom_array[33458] = 32'hFFFFFFF1;
    // rom_array[33459] = 32'hFFFFFFF1;
    // rom_array[33460] = 32'hFFFFFFF1;
    // rom_array[33461] = 32'hFFFFFFF1;
    // rom_array[33462] = 32'hFFFFFFF1;
    // rom_array[33463] = 32'hFFFFFFF1;
    // rom_array[33464] = 32'hFFFFFFF1;
    // rom_array[33465] = 32'hFFFFFFF0;
    // rom_array[33466] = 32'hFFFFFFF0;
    // rom_array[33467] = 32'hFFFFFFF1;
    // rom_array[33468] = 32'hFFFFFFF1;
    // rom_array[33469] = 32'hFFFFFFF0;
    // rom_array[33470] = 32'hFFFFFFF0;
    // rom_array[33471] = 32'hFFFFFFF1;
    // rom_array[33472] = 32'hFFFFFFF1;
    // rom_array[33473] = 32'hFFFFFFF0;
    // rom_array[33474] = 32'hFFFFFFF0;
    // rom_array[33475] = 32'hFFFFFFF1;
    // rom_array[33476] = 32'hFFFFFFF1;
    // rom_array[33477] = 32'hFFFFFFF0;
    // rom_array[33478] = 32'hFFFFFFF0;
    // rom_array[33479] = 32'hFFFFFFF1;
    // rom_array[33480] = 32'hFFFFFFF1;
    // rom_array[33481] = 32'hFFFFFFF0;
    // rom_array[33482] = 32'hFFFFFFF0;
    // rom_array[33483] = 32'hFFFFFFF1;
    // rom_array[33484] = 32'hFFFFFFF1;
    // rom_array[33485] = 32'hFFFFFFF0;
    // rom_array[33486] = 32'hFFFFFFF0;
    // rom_array[33487] = 32'hFFFFFFF1;
    // rom_array[33488] = 32'hFFFFFFF1;
    // rom_array[33489] = 32'hFFFFFFF0;
    // rom_array[33490] = 32'hFFFFFFF0;
    // rom_array[33491] = 32'hFFFFFFF1;
    // rom_array[33492] = 32'hFFFFFFF1;
    // rom_array[33493] = 32'hFFFFFFF0;
    // rom_array[33494] = 32'hFFFFFFF0;
    // rom_array[33495] = 32'hFFFFFFF1;
    // rom_array[33496] = 32'hFFFFFFF1;
    // rom_array[33497] = 32'hFFFFFFF1;
    // rom_array[33498] = 32'hFFFFFFF1;
    // rom_array[33499] = 32'hFFFFFFF1;
    // rom_array[33500] = 32'hFFFFFFF1;
    // rom_array[33501] = 32'hFFFFFFF0;
    // rom_array[33502] = 32'hFFFFFFF0;
    // rom_array[33503] = 32'hFFFFFFF0;
    // rom_array[33504] = 32'hFFFFFFF0;
    // rom_array[33505] = 32'hFFFFFFF1;
    // rom_array[33506] = 32'hFFFFFFF1;
    // rom_array[33507] = 32'hFFFFFFF1;
    // rom_array[33508] = 32'hFFFFFFF1;
    // rom_array[33509] = 32'hFFFFFFF0;
    // rom_array[33510] = 32'hFFFFFFF0;
    // rom_array[33511] = 32'hFFFFFFF0;
    // rom_array[33512] = 32'hFFFFFFF0;
    // rom_array[33513] = 32'hFFFFFFF1;
    // rom_array[33514] = 32'hFFFFFFF1;
    // rom_array[33515] = 32'hFFFFFFF1;
    // rom_array[33516] = 32'hFFFFFFF1;
    // rom_array[33517] = 32'hFFFFFFF1;
    // rom_array[33518] = 32'hFFFFFFF1;
    // rom_array[33519] = 32'hFFFFFFF1;
    // rom_array[33520] = 32'hFFFFFFF1;
    // rom_array[33521] = 32'hFFFFFFF1;
    // rom_array[33522] = 32'hFFFFFFF1;
    // rom_array[33523] = 32'hFFFFFFF1;
    // rom_array[33524] = 32'hFFFFFFF1;
    // rom_array[33525] = 32'hFFFFFFF1;
    // rom_array[33526] = 32'hFFFFFFF1;
    // rom_array[33527] = 32'hFFFFFFF1;
    // rom_array[33528] = 32'hFFFFFFF1;
    // rom_array[33529] = 32'hFFFFFFF1;
    // rom_array[33530] = 32'hFFFFFFF1;
    // rom_array[33531] = 32'hFFFFFFF1;
    // rom_array[33532] = 32'hFFFFFFF1;
    // rom_array[33533] = 32'hFFFFFFF1;
    // rom_array[33534] = 32'hFFFFFFF1;
    // rom_array[33535] = 32'hFFFFFFF0;
    // rom_array[33536] = 32'hFFFFFFF0;
    // rom_array[33537] = 32'hFFFFFFF1;
    // rom_array[33538] = 32'hFFFFFFF1;
    // rom_array[33539] = 32'hFFFFFFF1;
    // rom_array[33540] = 32'hFFFFFFF1;
    // rom_array[33541] = 32'hFFFFFFF1;
    // rom_array[33542] = 32'hFFFFFFF1;
    // rom_array[33543] = 32'hFFFFFFF0;
    // rom_array[33544] = 32'hFFFFFFF0;
    // rom_array[33545] = 32'hFFFFFFF0;
    // rom_array[33546] = 32'hFFFFFFF0;
    // rom_array[33547] = 32'hFFFFFFF1;
    // rom_array[33548] = 32'hFFFFFFF1;
    // rom_array[33549] = 32'hFFFFFFF0;
    // rom_array[33550] = 32'hFFFFFFF0;
    // rom_array[33551] = 32'hFFFFFFF0;
    // rom_array[33552] = 32'hFFFFFFF0;
    // rom_array[33553] = 32'hFFFFFFF0;
    // rom_array[33554] = 32'hFFFFFFF0;
    // rom_array[33555] = 32'hFFFFFFF1;
    // rom_array[33556] = 32'hFFFFFFF1;
    // rom_array[33557] = 32'hFFFFFFF0;
    // rom_array[33558] = 32'hFFFFFFF0;
    // rom_array[33559] = 32'hFFFFFFF0;
    // rom_array[33560] = 32'hFFFFFFF0;
    // rom_array[33561] = 32'hFFFFFFF1;
    // rom_array[33562] = 32'hFFFFFFF1;
    // rom_array[33563] = 32'hFFFFFFF1;
    // rom_array[33564] = 32'hFFFFFFF1;
    // rom_array[33565] = 32'hFFFFFFF0;
    // rom_array[33566] = 32'hFFFFFFF0;
    // rom_array[33567] = 32'hFFFFFFF0;
    // rom_array[33568] = 32'hFFFFFFF0;
    // rom_array[33569] = 32'hFFFFFFF1;
    // rom_array[33570] = 32'hFFFFFFF1;
    // rom_array[33571] = 32'hFFFFFFF1;
    // rom_array[33572] = 32'hFFFFFFF1;
    // rom_array[33573] = 32'hFFFFFFF0;
    // rom_array[33574] = 32'hFFFFFFF0;
    // rom_array[33575] = 32'hFFFFFFF0;
    // rom_array[33576] = 32'hFFFFFFF0;
    // rom_array[33577] = 32'hFFFFFFF1;
    // rom_array[33578] = 32'hFFFFFFF1;
    // rom_array[33579] = 32'hFFFFFFF1;
    // rom_array[33580] = 32'hFFFFFFF1;
    // rom_array[33581] = 32'hFFFFFFF0;
    // rom_array[33582] = 32'hFFFFFFF0;
    // rom_array[33583] = 32'hFFFFFFF0;
    // rom_array[33584] = 32'hFFFFFFF0;
    // rom_array[33585] = 32'hFFFFFFF1;
    // rom_array[33586] = 32'hFFFFFFF1;
    // rom_array[33587] = 32'hFFFFFFF1;
    // rom_array[33588] = 32'hFFFFFFF1;
    // rom_array[33589] = 32'hFFFFFFF0;
    // rom_array[33590] = 32'hFFFFFFF0;
    // rom_array[33591] = 32'hFFFFFFF0;
    // rom_array[33592] = 32'hFFFFFFF0;
    // rom_array[33593] = 32'hFFFFFFF1;
    // rom_array[33594] = 32'hFFFFFFF1;
    // rom_array[33595] = 32'hFFFFFFF1;
    // rom_array[33596] = 32'hFFFFFFF1;
    // rom_array[33597] = 32'hFFFFFFF0;
    // rom_array[33598] = 32'hFFFFFFF0;
    // rom_array[33599] = 32'hFFFFFFF0;
    // rom_array[33600] = 32'hFFFFFFF0;
    // rom_array[33601] = 32'hFFFFFFF1;
    // rom_array[33602] = 32'hFFFFFFF1;
    // rom_array[33603] = 32'hFFFFFFF1;
    // rom_array[33604] = 32'hFFFFFFF1;
    // rom_array[33605] = 32'hFFFFFFF0;
    // rom_array[33606] = 32'hFFFFFFF0;
    // rom_array[33607] = 32'hFFFFFFF0;
    // rom_array[33608] = 32'hFFFFFFF0;
    // rom_array[33609] = 32'hFFFFFFF1;
    // rom_array[33610] = 32'hFFFFFFF1;
    // rom_array[33611] = 32'hFFFFFFF1;
    // rom_array[33612] = 32'hFFFFFFF1;
    // rom_array[33613] = 32'hFFFFFFF0;
    // rom_array[33614] = 32'hFFFFFFF0;
    // rom_array[33615] = 32'hFFFFFFF0;
    // rom_array[33616] = 32'hFFFFFFF0;
    // rom_array[33617] = 32'hFFFFFFF1;
    // rom_array[33618] = 32'hFFFFFFF1;
    // rom_array[33619] = 32'hFFFFFFF1;
    // rom_array[33620] = 32'hFFFFFFF1;
    // rom_array[33621] = 32'hFFFFFFF0;
    // rom_array[33622] = 32'hFFFFFFF0;
    // rom_array[33623] = 32'hFFFFFFF0;
    // rom_array[33624] = 32'hFFFFFFF0;
    // rom_array[33625] = 32'hFFFFFFF1;
    // rom_array[33626] = 32'hFFFFFFF1;
    // rom_array[33627] = 32'hFFFFFFF1;
    // rom_array[33628] = 32'hFFFFFFF1;
    // rom_array[33629] = 32'hFFFFFFF0;
    // rom_array[33630] = 32'hFFFFFFF0;
    // rom_array[33631] = 32'hFFFFFFF0;
    // rom_array[33632] = 32'hFFFFFFF0;
    // rom_array[33633] = 32'hFFFFFFF1;
    // rom_array[33634] = 32'hFFFFFFF1;
    // rom_array[33635] = 32'hFFFFFFF1;
    // rom_array[33636] = 32'hFFFFFFF1;
    // rom_array[33637] = 32'hFFFFFFF0;
    // rom_array[33638] = 32'hFFFFFFF0;
    // rom_array[33639] = 32'hFFFFFFF0;
    // rom_array[33640] = 32'hFFFFFFF0;
    // rom_array[33641] = 32'hFFFFFFF1;
    // rom_array[33642] = 32'hFFFFFFF1;
    // rom_array[33643] = 32'hFFFFFFF1;
    // rom_array[33644] = 32'hFFFFFFF1;
    // rom_array[33645] = 32'hFFFFFFF0;
    // rom_array[33646] = 32'hFFFFFFF0;
    // rom_array[33647] = 32'hFFFFFFF0;
    // rom_array[33648] = 32'hFFFFFFF0;
    // rom_array[33649] = 32'hFFFFFFF1;
    // rom_array[33650] = 32'hFFFFFFF1;
    // rom_array[33651] = 32'hFFFFFFF1;
    // rom_array[33652] = 32'hFFFFFFF1;
    // rom_array[33653] = 32'hFFFFFFF0;
    // rom_array[33654] = 32'hFFFFFFF0;
    // rom_array[33655] = 32'hFFFFFFF0;
    // rom_array[33656] = 32'hFFFFFFF0;
    // rom_array[33657] = 32'hFFFFFFF1;
    // rom_array[33658] = 32'hFFFFFFF1;
    // rom_array[33659] = 32'hFFFFFFF1;
    // rom_array[33660] = 32'hFFFFFFF1;
    // rom_array[33661] = 32'hFFFFFFF0;
    // rom_array[33662] = 32'hFFFFFFF0;
    // rom_array[33663] = 32'hFFFFFFF0;
    // rom_array[33664] = 32'hFFFFFFF0;
    // rom_array[33665] = 32'hFFFFFFF1;
    // rom_array[33666] = 32'hFFFFFFF1;
    // rom_array[33667] = 32'hFFFFFFF1;
    // rom_array[33668] = 32'hFFFFFFF1;
    // rom_array[33669] = 32'hFFFFFFF0;
    // rom_array[33670] = 32'hFFFFFFF0;
    // rom_array[33671] = 32'hFFFFFFF0;
    // rom_array[33672] = 32'hFFFFFFF0;
    // rom_array[33673] = 32'hFFFFFFF1;
    // rom_array[33674] = 32'hFFFFFFF1;
    // rom_array[33675] = 32'hFFFFFFF1;
    // rom_array[33676] = 32'hFFFFFFF1;
    // rom_array[33677] = 32'hFFFFFFF0;
    // rom_array[33678] = 32'hFFFFFFF0;
    // rom_array[33679] = 32'hFFFFFFF0;
    // rom_array[33680] = 32'hFFFFFFF0;
    // rom_array[33681] = 32'hFFFFFFF1;
    // rom_array[33682] = 32'hFFFFFFF1;
    // rom_array[33683] = 32'hFFFFFFF1;
    // rom_array[33684] = 32'hFFFFFFF1;
    // rom_array[33685] = 32'hFFFFFFF0;
    // rom_array[33686] = 32'hFFFFFFF0;
    // rom_array[33687] = 32'hFFFFFFF0;
    // rom_array[33688] = 32'hFFFFFFF0;
    // rom_array[33689] = 32'hFFFFFFF1;
    // rom_array[33690] = 32'hFFFFFFF1;
    // rom_array[33691] = 32'hFFFFFFF1;
    // rom_array[33692] = 32'hFFFFFFF1;
    // rom_array[33693] = 32'hFFFFFFF0;
    // rom_array[33694] = 32'hFFFFFFF0;
    // rom_array[33695] = 32'hFFFFFFF0;
    // rom_array[33696] = 32'hFFFFFFF0;
    // rom_array[33697] = 32'hFFFFFFF1;
    // rom_array[33698] = 32'hFFFFFFF1;
    // rom_array[33699] = 32'hFFFFFFF1;
    // rom_array[33700] = 32'hFFFFFFF1;
    // rom_array[33701] = 32'hFFFFFFF0;
    // rom_array[33702] = 32'hFFFFFFF0;
    // rom_array[33703] = 32'hFFFFFFF0;
    // rom_array[33704] = 32'hFFFFFFF0;
    // rom_array[33705] = 32'hFFFFFFF1;
    // rom_array[33706] = 32'hFFFFFFF1;
    // rom_array[33707] = 32'hFFFFFFF1;
    // rom_array[33708] = 32'hFFFFFFF1;
    // rom_array[33709] = 32'hFFFFFFF0;
    // rom_array[33710] = 32'hFFFFFFF0;
    // rom_array[33711] = 32'hFFFFFFF0;
    // rom_array[33712] = 32'hFFFFFFF0;
    // rom_array[33713] = 32'hFFFFFFF1;
    // rom_array[33714] = 32'hFFFFFFF1;
    // rom_array[33715] = 32'hFFFFFFF1;
    // rom_array[33716] = 32'hFFFFFFF1;
    // rom_array[33717] = 32'hFFFFFFF0;
    // rom_array[33718] = 32'hFFFFFFF0;
    // rom_array[33719] = 32'hFFFFFFF0;
    // rom_array[33720] = 32'hFFFFFFF0;
    // rom_array[33721] = 32'hFFFFFFF1;
    // rom_array[33722] = 32'hFFFFFFF1;
    // rom_array[33723] = 32'hFFFFFFF1;
    // rom_array[33724] = 32'hFFFFFFF1;
    // rom_array[33725] = 32'hFFFFFFF0;
    // rom_array[33726] = 32'hFFFFFFF0;
    // rom_array[33727] = 32'hFFFFFFF0;
    // rom_array[33728] = 32'hFFFFFFF0;
    // rom_array[33729] = 32'hFFFFFFF1;
    // rom_array[33730] = 32'hFFFFFFF1;
    // rom_array[33731] = 32'hFFFFFFF1;
    // rom_array[33732] = 32'hFFFFFFF1;
    // rom_array[33733] = 32'hFFFFFFF0;
    // rom_array[33734] = 32'hFFFFFFF0;
    // rom_array[33735] = 32'hFFFFFFF0;
    // rom_array[33736] = 32'hFFFFFFF0;
    // rom_array[33737] = 32'hFFFFFFF0;
    // rom_array[33738] = 32'hFFFFFFF0;
    // rom_array[33739] = 32'hFFFFFFF0;
    // rom_array[33740] = 32'hFFFFFFF0;
    // rom_array[33741] = 32'hFFFFFFF0;
    // rom_array[33742] = 32'hFFFFFFF0;
    // rom_array[33743] = 32'hFFFFFFF1;
    // rom_array[33744] = 32'hFFFFFFF1;
    // rom_array[33745] = 32'hFFFFFFF0;
    // rom_array[33746] = 32'hFFFFFFF0;
    // rom_array[33747] = 32'hFFFFFFF0;
    // rom_array[33748] = 32'hFFFFFFF0;
    // rom_array[33749] = 32'hFFFFFFF0;
    // rom_array[33750] = 32'hFFFFFFF0;
    // rom_array[33751] = 32'hFFFFFFF1;
    // rom_array[33752] = 32'hFFFFFFF1;
    // rom_array[33753] = 32'hFFFFFFF0;
    // rom_array[33754] = 32'hFFFFFFF0;
    // rom_array[33755] = 32'hFFFFFFF0;
    // rom_array[33756] = 32'hFFFFFFF0;
    // rom_array[33757] = 32'hFFFFFFF1;
    // rom_array[33758] = 32'hFFFFFFF1;
    // rom_array[33759] = 32'hFFFFFFF1;
    // rom_array[33760] = 32'hFFFFFFF1;
    // rom_array[33761] = 32'hFFFFFFF0;
    // rom_array[33762] = 32'hFFFFFFF0;
    // rom_array[33763] = 32'hFFFFFFF0;
    // rom_array[33764] = 32'hFFFFFFF0;
    // rom_array[33765] = 32'hFFFFFFF1;
    // rom_array[33766] = 32'hFFFFFFF1;
    // rom_array[33767] = 32'hFFFFFFF1;
    // rom_array[33768] = 32'hFFFFFFF1;
    // rom_array[33769] = 32'hFFFFFFF0;
    // rom_array[33770] = 32'hFFFFFFF0;
    // rom_array[33771] = 32'hFFFFFFF1;
    // rom_array[33772] = 32'hFFFFFFF1;
    // rom_array[33773] = 32'hFFFFFFF0;
    // rom_array[33774] = 32'hFFFFFFF0;
    // rom_array[33775] = 32'hFFFFFFF1;
    // rom_array[33776] = 32'hFFFFFFF1;
    // rom_array[33777] = 32'hFFFFFFF0;
    // rom_array[33778] = 32'hFFFFFFF0;
    // rom_array[33779] = 32'hFFFFFFF1;
    // rom_array[33780] = 32'hFFFFFFF1;
    // rom_array[33781] = 32'hFFFFFFF0;
    // rom_array[33782] = 32'hFFFFFFF0;
    // rom_array[33783] = 32'hFFFFFFF1;
    // rom_array[33784] = 32'hFFFFFFF1;
    // rom_array[33785] = 32'hFFFFFFF0;
    // rom_array[33786] = 32'hFFFFFFF0;
    // rom_array[33787] = 32'hFFFFFFF0;
    // rom_array[33788] = 32'hFFFFFFF0;
    // rom_array[33789] = 32'hFFFFFFF1;
    // rom_array[33790] = 32'hFFFFFFF1;
    // rom_array[33791] = 32'hFFFFFFF1;
    // rom_array[33792] = 32'hFFFFFFF1;
    // rom_array[33793] = 32'hFFFFFFF0;
    // rom_array[33794] = 32'hFFFFFFF0;
    // rom_array[33795] = 32'hFFFFFFF0;
    // rom_array[33796] = 32'hFFFFFFF0;
    // rom_array[33797] = 32'hFFFFFFF1;
    // rom_array[33798] = 32'hFFFFFFF1;
    // rom_array[33799] = 32'hFFFFFFF1;
    // rom_array[33800] = 32'hFFFFFFF1;
    // rom_array[33801] = 32'hFFFFFFF0;
    // rom_array[33802] = 32'hFFFFFFF0;
    // rom_array[33803] = 32'hFFFFFFF0;
    // rom_array[33804] = 32'hFFFFFFF0;
    // rom_array[33805] = 32'hFFFFFFF1;
    // rom_array[33806] = 32'hFFFFFFF1;
    // rom_array[33807] = 32'hFFFFFFF1;
    // rom_array[33808] = 32'hFFFFFFF1;
    // rom_array[33809] = 32'hFFFFFFF0;
    // rom_array[33810] = 32'hFFFFFFF0;
    // rom_array[33811] = 32'hFFFFFFF0;
    // rom_array[33812] = 32'hFFFFFFF0;
    // rom_array[33813] = 32'hFFFFFFF1;
    // rom_array[33814] = 32'hFFFFFFF1;
    // rom_array[33815] = 32'hFFFFFFF1;
    // rom_array[33816] = 32'hFFFFFFF1;
    // rom_array[33817] = 32'hFFFFFFF0;
    // rom_array[33818] = 32'hFFFFFFF0;
    // rom_array[33819] = 32'hFFFFFFF1;
    // rom_array[33820] = 32'hFFFFFFF1;
    // rom_array[33821] = 32'hFFFFFFF0;
    // rom_array[33822] = 32'hFFFFFFF0;
    // rom_array[33823] = 32'hFFFFFFF1;
    // rom_array[33824] = 32'hFFFFFFF1;
    // rom_array[33825] = 32'hFFFFFFF0;
    // rom_array[33826] = 32'hFFFFFFF0;
    // rom_array[33827] = 32'hFFFFFFF1;
    // rom_array[33828] = 32'hFFFFFFF1;
    // rom_array[33829] = 32'hFFFFFFF0;
    // rom_array[33830] = 32'hFFFFFFF0;
    // rom_array[33831] = 32'hFFFFFFF1;
    // rom_array[33832] = 32'hFFFFFFF1;
    // rom_array[33833] = 32'hFFFFFFF0;
    // rom_array[33834] = 32'hFFFFFFF0;
    // rom_array[33835] = 32'hFFFFFFF1;
    // rom_array[33836] = 32'hFFFFFFF1;
    // rom_array[33837] = 32'hFFFFFFF0;
    // rom_array[33838] = 32'hFFFFFFF0;
    // rom_array[33839] = 32'hFFFFFFF1;
    // rom_array[33840] = 32'hFFFFFFF1;
    // rom_array[33841] = 32'hFFFFFFF0;
    // rom_array[33842] = 32'hFFFFFFF0;
    // rom_array[33843] = 32'hFFFFFFF1;
    // rom_array[33844] = 32'hFFFFFFF1;
    // rom_array[33845] = 32'hFFFFFFF0;
    // rom_array[33846] = 32'hFFFFFFF0;
    // rom_array[33847] = 32'hFFFFFFF1;
    // rom_array[33848] = 32'hFFFFFFF1;
    // rom_array[33849] = 32'hFFFFFFF0;
    // rom_array[33850] = 32'hFFFFFFF0;
    // rom_array[33851] = 32'hFFFFFFF0;
    // rom_array[33852] = 32'hFFFFFFF0;
    // rom_array[33853] = 32'hFFFFFFF1;
    // rom_array[33854] = 32'hFFFFFFF1;
    // rom_array[33855] = 32'hFFFFFFF1;
    // rom_array[33856] = 32'hFFFFFFF1;
    // rom_array[33857] = 32'hFFFFFFF0;
    // rom_array[33858] = 32'hFFFFFFF0;
    // rom_array[33859] = 32'hFFFFFFF0;
    // rom_array[33860] = 32'hFFFFFFF0;
    // rom_array[33861] = 32'hFFFFFFF1;
    // rom_array[33862] = 32'hFFFFFFF1;
    // rom_array[33863] = 32'hFFFFFFF1;
    // rom_array[33864] = 32'hFFFFFFF1;
    // rom_array[33865] = 32'hFFFFFFF0;
    // rom_array[33866] = 32'hFFFFFFF0;
    // rom_array[33867] = 32'hFFFFFFF0;
    // rom_array[33868] = 32'hFFFFFFF0;
    // rom_array[33869] = 32'hFFFFFFF1;
    // rom_array[33870] = 32'hFFFFFFF1;
    // rom_array[33871] = 32'hFFFFFFF1;
    // rom_array[33872] = 32'hFFFFFFF1;
    // rom_array[33873] = 32'hFFFFFFF0;
    // rom_array[33874] = 32'hFFFFFFF0;
    // rom_array[33875] = 32'hFFFFFFF0;
    // rom_array[33876] = 32'hFFFFFFF0;
    // rom_array[33877] = 32'hFFFFFFF1;
    // rom_array[33878] = 32'hFFFFFFF1;
    // rom_array[33879] = 32'hFFFFFFF1;
    // rom_array[33880] = 32'hFFFFFFF1;
    // rom_array[33881] = 32'hFFFFFFF0;
    // rom_array[33882] = 32'hFFFFFFF0;
    // rom_array[33883] = 32'hFFFFFFF0;
    // rom_array[33884] = 32'hFFFFFFF0;
    // rom_array[33885] = 32'hFFFFFFF1;
    // rom_array[33886] = 32'hFFFFFFF1;
    // rom_array[33887] = 32'hFFFFFFF1;
    // rom_array[33888] = 32'hFFFFFFF1;
    // rom_array[33889] = 32'hFFFFFFF0;
    // rom_array[33890] = 32'hFFFFFFF0;
    // rom_array[33891] = 32'hFFFFFFF0;
    // rom_array[33892] = 32'hFFFFFFF0;
    // rom_array[33893] = 32'hFFFFFFF1;
    // rom_array[33894] = 32'hFFFFFFF1;
    // rom_array[33895] = 32'hFFFFFFF1;
    // rom_array[33896] = 32'hFFFFFFF1;
    // rom_array[33897] = 32'hFFFFFFF0;
    // rom_array[33898] = 32'hFFFFFFF0;
    // rom_array[33899] = 32'hFFFFFFF0;
    // rom_array[33900] = 32'hFFFFFFF0;
    // rom_array[33901] = 32'hFFFFFFF1;
    // rom_array[33902] = 32'hFFFFFFF1;
    // rom_array[33903] = 32'hFFFFFFF1;
    // rom_array[33904] = 32'hFFFFFFF1;
    // rom_array[33905] = 32'hFFFFFFF0;
    // rom_array[33906] = 32'hFFFFFFF0;
    // rom_array[33907] = 32'hFFFFFFF0;
    // rom_array[33908] = 32'hFFFFFFF0;
    // rom_array[33909] = 32'hFFFFFFF1;
    // rom_array[33910] = 32'hFFFFFFF1;
    // rom_array[33911] = 32'hFFFFFFF1;
    // rom_array[33912] = 32'hFFFFFFF1;
    // rom_array[33913] = 32'hFFFFFFF0;
    // rom_array[33914] = 32'hFFFFFFF0;
    // rom_array[33915] = 32'hFFFFFFF0;
    // rom_array[33916] = 32'hFFFFFFF0;
    // rom_array[33917] = 32'hFFFFFFF1;
    // rom_array[33918] = 32'hFFFFFFF1;
    // rom_array[33919] = 32'hFFFFFFF1;
    // rom_array[33920] = 32'hFFFFFFF1;
    // rom_array[33921] = 32'hFFFFFFF0;
    // rom_array[33922] = 32'hFFFFFFF0;
    // rom_array[33923] = 32'hFFFFFFF0;
    // rom_array[33924] = 32'hFFFFFFF0;
    // rom_array[33925] = 32'hFFFFFFF1;
    // rom_array[33926] = 32'hFFFFFFF1;
    // rom_array[33927] = 32'hFFFFFFF1;
    // rom_array[33928] = 32'hFFFFFFF1;
    // rom_array[33929] = 32'hFFFFFFF0;
    // rom_array[33930] = 32'hFFFFFFF0;
    // rom_array[33931] = 32'hFFFFFFF0;
    // rom_array[33932] = 32'hFFFFFFF0;
    // rom_array[33933] = 32'hFFFFFFF1;
    // rom_array[33934] = 32'hFFFFFFF1;
    // rom_array[33935] = 32'hFFFFFFF1;
    // rom_array[33936] = 32'hFFFFFFF1;
    // rom_array[33937] = 32'hFFFFFFF0;
    // rom_array[33938] = 32'hFFFFFFF0;
    // rom_array[33939] = 32'hFFFFFFF0;
    // rom_array[33940] = 32'hFFFFFFF0;
    // rom_array[33941] = 32'hFFFFFFF1;
    // rom_array[33942] = 32'hFFFFFFF1;
    // rom_array[33943] = 32'hFFFFFFF1;
    // rom_array[33944] = 32'hFFFFFFF1;
    // rom_array[33945] = 32'hFFFFFFF0;
    // rom_array[33946] = 32'hFFFFFFF0;
    // rom_array[33947] = 32'hFFFFFFF0;
    // rom_array[33948] = 32'hFFFFFFF0;
    // rom_array[33949] = 32'hFFFFFFF1;
    // rom_array[33950] = 32'hFFFFFFF1;
    // rom_array[33951] = 32'hFFFFFFF1;
    // rom_array[33952] = 32'hFFFFFFF1;
    // rom_array[33953] = 32'hFFFFFFF0;
    // rom_array[33954] = 32'hFFFFFFF0;
    // rom_array[33955] = 32'hFFFFFFF0;
    // rom_array[33956] = 32'hFFFFFFF0;
    // rom_array[33957] = 32'hFFFFFFF1;
    // rom_array[33958] = 32'hFFFFFFF1;
    // rom_array[33959] = 32'hFFFFFFF1;
    // rom_array[33960] = 32'hFFFFFFF1;
    // rom_array[33961] = 32'hFFFFFFF0;
    // rom_array[33962] = 32'hFFFFFFF0;
    // rom_array[33963] = 32'hFFFFFFF0;
    // rom_array[33964] = 32'hFFFFFFF0;
    // rom_array[33965] = 32'hFFFFFFF1;
    // rom_array[33966] = 32'hFFFFFFF1;
    // rom_array[33967] = 32'hFFFFFFF1;
    // rom_array[33968] = 32'hFFFFFFF1;
    // rom_array[33969] = 32'hFFFFFFF0;
    // rom_array[33970] = 32'hFFFFFFF0;
    // rom_array[33971] = 32'hFFFFFFF0;
    // rom_array[33972] = 32'hFFFFFFF0;
    // rom_array[33973] = 32'hFFFFFFF1;
    // rom_array[33974] = 32'hFFFFFFF1;
    // rom_array[33975] = 32'hFFFFFFF1;
    // rom_array[33976] = 32'hFFFFFFF1;
    // rom_array[33977] = 32'hFFFFFFF0;
    // rom_array[33978] = 32'hFFFFFFF0;
    // rom_array[33979] = 32'hFFFFFFF1;
    // rom_array[33980] = 32'hFFFFFFF1;
    // rom_array[33981] = 32'hFFFFFFF0;
    // rom_array[33982] = 32'hFFFFFFF0;
    // rom_array[33983] = 32'hFFFFFFF1;
    // rom_array[33984] = 32'hFFFFFFF1;
    // rom_array[33985] = 32'hFFFFFFF0;
    // rom_array[33986] = 32'hFFFFFFF0;
    // rom_array[33987] = 32'hFFFFFFF1;
    // rom_array[33988] = 32'hFFFFFFF1;
    // rom_array[33989] = 32'hFFFFFFF0;
    // rom_array[33990] = 32'hFFFFFFF0;
    // rom_array[33991] = 32'hFFFFFFF1;
    // rom_array[33992] = 32'hFFFFFFF1;
    // rom_array[33993] = 32'hFFFFFFF1;
    // rom_array[33994] = 32'hFFFFFFF1;
    // rom_array[33995] = 32'hFFFFFFF1;
    // rom_array[33996] = 32'hFFFFFFF1;
    // rom_array[33997] = 32'hFFFFFFF1;
    // rom_array[33998] = 32'hFFFFFFF1;
    // rom_array[33999] = 32'hFFFFFFF1;
    // rom_array[34000] = 32'hFFFFFFF1;
    // rom_array[34001] = 32'hFFFFFFF1;
    // rom_array[34002] = 32'hFFFFFFF1;
    // rom_array[34003] = 32'hFFFFFFF1;
    // rom_array[34004] = 32'hFFFFFFF1;
    // rom_array[34005] = 32'hFFFFFFF1;
    // rom_array[34006] = 32'hFFFFFFF1;
    // rom_array[34007] = 32'hFFFFFFF1;
    // rom_array[34008] = 32'hFFFFFFF1;
    // rom_array[34009] = 32'hFFFFFFF0;
    // rom_array[34010] = 32'hFFFFFFF0;
    // rom_array[34011] = 32'hFFFFFFF1;
    // rom_array[34012] = 32'hFFFFFFF1;
    // rom_array[34013] = 32'hFFFFFFF0;
    // rom_array[34014] = 32'hFFFFFFF0;
    // rom_array[34015] = 32'hFFFFFFF1;
    // rom_array[34016] = 32'hFFFFFFF1;
    // rom_array[34017] = 32'hFFFFFFF0;
    // rom_array[34018] = 32'hFFFFFFF0;
    // rom_array[34019] = 32'hFFFFFFF1;
    // rom_array[34020] = 32'hFFFFFFF1;
    // rom_array[34021] = 32'hFFFFFFF0;
    // rom_array[34022] = 32'hFFFFFFF0;
    // rom_array[34023] = 32'hFFFFFFF1;
    // rom_array[34024] = 32'hFFFFFFF1;
    // rom_array[34025] = 32'hFFFFFFF1;
    // rom_array[34026] = 32'hFFFFFFF1;
    // rom_array[34027] = 32'hFFFFFFF1;
    // rom_array[34028] = 32'hFFFFFFF1;
    // rom_array[34029] = 32'hFFFFFFF1;
    // rom_array[34030] = 32'hFFFFFFF1;
    // rom_array[34031] = 32'hFFFFFFF1;
    // rom_array[34032] = 32'hFFFFFFF1;
    // rom_array[34033] = 32'hFFFFFFF1;
    // rom_array[34034] = 32'hFFFFFFF1;
    // rom_array[34035] = 32'hFFFFFFF1;
    // rom_array[34036] = 32'hFFFFFFF1;
    // rom_array[34037] = 32'hFFFFFFF1;
    // rom_array[34038] = 32'hFFFFFFF1;
    // rom_array[34039] = 32'hFFFFFFF1;
    // rom_array[34040] = 32'hFFFFFFF1;
    // rom_array[34041] = 32'hFFFFFFF1;
    // rom_array[34042] = 32'hFFFFFFF1;
    // rom_array[34043] = 32'hFFFFFFF1;
    // rom_array[34044] = 32'hFFFFFFF1;
    // rom_array[34045] = 32'hFFFFFFF1;
    // rom_array[34046] = 32'hFFFFFFF1;
    // rom_array[34047] = 32'hFFFFFFF1;
    // rom_array[34048] = 32'hFFFFFFF1;
    // rom_array[34049] = 32'hFFFFFFF1;
    // rom_array[34050] = 32'hFFFFFFF1;
    // rom_array[34051] = 32'hFFFFFFF1;
    // rom_array[34052] = 32'hFFFFFFF1;
    // rom_array[34053] = 32'hFFFFFFF1;
    // rom_array[34054] = 32'hFFFFFFF1;
    // rom_array[34055] = 32'hFFFFFFF1;
    // rom_array[34056] = 32'hFFFFFFF1;
    // rom_array[34057] = 32'hFFFFFFF0;
    // rom_array[34058] = 32'hFFFFFFF0;
    // rom_array[34059] = 32'hFFFFFFF1;
    // rom_array[34060] = 32'hFFFFFFF1;
    // rom_array[34061] = 32'hFFFFFFF0;
    // rom_array[34062] = 32'hFFFFFFF0;
    // rom_array[34063] = 32'hFFFFFFF1;
    // rom_array[34064] = 32'hFFFFFFF1;
    // rom_array[34065] = 32'hFFFFFFF0;
    // rom_array[34066] = 32'hFFFFFFF0;
    // rom_array[34067] = 32'hFFFFFFF1;
    // rom_array[34068] = 32'hFFFFFFF1;
    // rom_array[34069] = 32'hFFFFFFF0;
    // rom_array[34070] = 32'hFFFFFFF0;
    // rom_array[34071] = 32'hFFFFFFF1;
    // rom_array[34072] = 32'hFFFFFFF1;
    // rom_array[34073] = 32'hFFFFFFF0;
    // rom_array[34074] = 32'hFFFFFFF0;
    // rom_array[34075] = 32'hFFFFFFF1;
    // rom_array[34076] = 32'hFFFFFFF1;
    // rom_array[34077] = 32'hFFFFFFF0;
    // rom_array[34078] = 32'hFFFFFFF0;
    // rom_array[34079] = 32'hFFFFFFF1;
    // rom_array[34080] = 32'hFFFFFFF1;
    // rom_array[34081] = 32'hFFFFFFF0;
    // rom_array[34082] = 32'hFFFFFFF0;
    // rom_array[34083] = 32'hFFFFFFF1;
    // rom_array[34084] = 32'hFFFFFFF1;
    // rom_array[34085] = 32'hFFFFFFF0;
    // rom_array[34086] = 32'hFFFFFFF0;
    // rom_array[34087] = 32'hFFFFFFF1;
    // rom_array[34088] = 32'hFFFFFFF1;
    // rom_array[34089] = 32'hFFFFFFF0;
    // rom_array[34090] = 32'hFFFFFFF0;
    // rom_array[34091] = 32'hFFFFFFF1;
    // rom_array[34092] = 32'hFFFFFFF1;
    // rom_array[34093] = 32'hFFFFFFF0;
    // rom_array[34094] = 32'hFFFFFFF0;
    // rom_array[34095] = 32'hFFFFFFF1;
    // rom_array[34096] = 32'hFFFFFFF1;
    // rom_array[34097] = 32'hFFFFFFF0;
    // rom_array[34098] = 32'hFFFFFFF0;
    // rom_array[34099] = 32'hFFFFFFF1;
    // rom_array[34100] = 32'hFFFFFFF1;
    // rom_array[34101] = 32'hFFFFFFF0;
    // rom_array[34102] = 32'hFFFFFFF0;
    // rom_array[34103] = 32'hFFFFFFF1;
    // rom_array[34104] = 32'hFFFFFFF1;
    // rom_array[34105] = 32'hFFFFFFF0;
    // rom_array[34106] = 32'hFFFFFFF0;
    // rom_array[34107] = 32'hFFFFFFF1;
    // rom_array[34108] = 32'hFFFFFFF1;
    // rom_array[34109] = 32'hFFFFFFF0;
    // rom_array[34110] = 32'hFFFFFFF0;
    // rom_array[34111] = 32'hFFFFFFF1;
    // rom_array[34112] = 32'hFFFFFFF1;
    // rom_array[34113] = 32'hFFFFFFF0;
    // rom_array[34114] = 32'hFFFFFFF0;
    // rom_array[34115] = 32'hFFFFFFF1;
    // rom_array[34116] = 32'hFFFFFFF1;
    // rom_array[34117] = 32'hFFFFFFF0;
    // rom_array[34118] = 32'hFFFFFFF0;
    // rom_array[34119] = 32'hFFFFFFF1;
    // rom_array[34120] = 32'hFFFFFFF1;
    // rom_array[34121] = 32'hFFFFFFF0;
    // rom_array[34122] = 32'hFFFFFFF0;
    // rom_array[34123] = 32'hFFFFFFF1;
    // rom_array[34124] = 32'hFFFFFFF1;
    // rom_array[34125] = 32'hFFFFFFF0;
    // rom_array[34126] = 32'hFFFFFFF0;
    // rom_array[34127] = 32'hFFFFFFF1;
    // rom_array[34128] = 32'hFFFFFFF1;
    // rom_array[34129] = 32'hFFFFFFF0;
    // rom_array[34130] = 32'hFFFFFFF0;
    // rom_array[34131] = 32'hFFFFFFF1;
    // rom_array[34132] = 32'hFFFFFFF1;
    // rom_array[34133] = 32'hFFFFFFF0;
    // rom_array[34134] = 32'hFFFFFFF0;
    // rom_array[34135] = 32'hFFFFFFF1;
    // rom_array[34136] = 32'hFFFFFFF1;
    // rom_array[34137] = 32'hFFFFFFF0;
    // rom_array[34138] = 32'hFFFFFFF0;
    // rom_array[34139] = 32'hFFFFFFF1;
    // rom_array[34140] = 32'hFFFFFFF1;
    // rom_array[34141] = 32'hFFFFFFF0;
    // rom_array[34142] = 32'hFFFFFFF0;
    // rom_array[34143] = 32'hFFFFFFF1;
    // rom_array[34144] = 32'hFFFFFFF1;
    // rom_array[34145] = 32'hFFFFFFF0;
    // rom_array[34146] = 32'hFFFFFFF0;
    // rom_array[34147] = 32'hFFFFFFF1;
    // rom_array[34148] = 32'hFFFFFFF1;
    // rom_array[34149] = 32'hFFFFFFF0;
    // rom_array[34150] = 32'hFFFFFFF0;
    // rom_array[34151] = 32'hFFFFFFF1;
    // rom_array[34152] = 32'hFFFFFFF1;
    // rom_array[34153] = 32'hFFFFFFF1;
    // rom_array[34154] = 32'hFFFFFFF1;
    // rom_array[34155] = 32'hFFFFFFF1;
    // rom_array[34156] = 32'hFFFFFFF1;
    // rom_array[34157] = 32'hFFFFFFF1;
    // rom_array[34158] = 32'hFFFFFFF1;
    // rom_array[34159] = 32'hFFFFFFF1;
    // rom_array[34160] = 32'hFFFFFFF1;
    // rom_array[34161] = 32'hFFFFFFF1;
    // rom_array[34162] = 32'hFFFFFFF1;
    // rom_array[34163] = 32'hFFFFFFF1;
    // rom_array[34164] = 32'hFFFFFFF1;
    // rom_array[34165] = 32'hFFFFFFF1;
    // rom_array[34166] = 32'hFFFFFFF1;
    // rom_array[34167] = 32'hFFFFFFF1;
    // rom_array[34168] = 32'hFFFFFFF1;
    // rom_array[34169] = 32'hFFFFFFF1;
    // rom_array[34170] = 32'hFFFFFFF1;
    // rom_array[34171] = 32'hFFFFFFF1;
    // rom_array[34172] = 32'hFFFFFFF1;
    // rom_array[34173] = 32'hFFFFFFF0;
    // rom_array[34174] = 32'hFFFFFFF0;
    // rom_array[34175] = 32'hFFFFFFF0;
    // rom_array[34176] = 32'hFFFFFFF0;
    // rom_array[34177] = 32'hFFFFFFF1;
    // rom_array[34178] = 32'hFFFFFFF1;
    // rom_array[34179] = 32'hFFFFFFF1;
    // rom_array[34180] = 32'hFFFFFFF1;
    // rom_array[34181] = 32'hFFFFFFF0;
    // rom_array[34182] = 32'hFFFFFFF0;
    // rom_array[34183] = 32'hFFFFFFF0;
    // rom_array[34184] = 32'hFFFFFFF0;
    // rom_array[34185] = 32'hFFFFFFF1;
    // rom_array[34186] = 32'hFFFFFFF1;
    // rom_array[34187] = 32'hFFFFFFF1;
    // rom_array[34188] = 32'hFFFFFFF1;
    // rom_array[34189] = 32'hFFFFFFF1;
    // rom_array[34190] = 32'hFFFFFFF1;
    // rom_array[34191] = 32'hFFFFFFF1;
    // rom_array[34192] = 32'hFFFFFFF1;
    // rom_array[34193] = 32'hFFFFFFF1;
    // rom_array[34194] = 32'hFFFFFFF1;
    // rom_array[34195] = 32'hFFFFFFF1;
    // rom_array[34196] = 32'hFFFFFFF1;
    // rom_array[34197] = 32'hFFFFFFF1;
    // rom_array[34198] = 32'hFFFFFFF1;
    // rom_array[34199] = 32'hFFFFFFF1;
    // rom_array[34200] = 32'hFFFFFFF1;
    // rom_array[34201] = 32'hFFFFFFF1;
    // rom_array[34202] = 32'hFFFFFFF1;
    // rom_array[34203] = 32'hFFFFFFF1;
    // rom_array[34204] = 32'hFFFFFFF1;
    // rom_array[34205] = 32'hFFFFFFF0;
    // rom_array[34206] = 32'hFFFFFFF0;
    // rom_array[34207] = 32'hFFFFFFF0;
    // rom_array[34208] = 32'hFFFFFFF0;
    // rom_array[34209] = 32'hFFFFFFF1;
    // rom_array[34210] = 32'hFFFFFFF1;
    // rom_array[34211] = 32'hFFFFFFF1;
    // rom_array[34212] = 32'hFFFFFFF1;
    // rom_array[34213] = 32'hFFFFFFF0;
    // rom_array[34214] = 32'hFFFFFFF0;
    // rom_array[34215] = 32'hFFFFFFF0;
    // rom_array[34216] = 32'hFFFFFFF0;
    // rom_array[34217] = 32'hFFFFFFF1;
    // rom_array[34218] = 32'hFFFFFFF1;
    // rom_array[34219] = 32'hFFFFFFF1;
    // rom_array[34220] = 32'hFFFFFFF1;
    // rom_array[34221] = 32'hFFFFFFF0;
    // rom_array[34222] = 32'hFFFFFFF0;
    // rom_array[34223] = 32'hFFFFFFF0;
    // rom_array[34224] = 32'hFFFFFFF0;
    // rom_array[34225] = 32'hFFFFFFF1;
    // rom_array[34226] = 32'hFFFFFFF1;
    // rom_array[34227] = 32'hFFFFFFF1;
    // rom_array[34228] = 32'hFFFFFFF1;
    // rom_array[34229] = 32'hFFFFFFF0;
    // rom_array[34230] = 32'hFFFFFFF0;
    // rom_array[34231] = 32'hFFFFFFF0;
    // rom_array[34232] = 32'hFFFFFFF0;
    // rom_array[34233] = 32'hFFFFFFF1;
    // rom_array[34234] = 32'hFFFFFFF1;
    // rom_array[34235] = 32'hFFFFFFF1;
    // rom_array[34236] = 32'hFFFFFFF1;
    // rom_array[34237] = 32'hFFFFFFF1;
    // rom_array[34238] = 32'hFFFFFFF1;
    // rom_array[34239] = 32'hFFFFFFF1;
    // rom_array[34240] = 32'hFFFFFFF1;
    // rom_array[34241] = 32'hFFFFFFF1;
    // rom_array[34242] = 32'hFFFFFFF1;
    // rom_array[34243] = 32'hFFFFFFF1;
    // rom_array[34244] = 32'hFFFFFFF1;
    // rom_array[34245] = 32'hFFFFFFF1;
    // rom_array[34246] = 32'hFFFFFFF1;
    // rom_array[34247] = 32'hFFFFFFF1;
    // rom_array[34248] = 32'hFFFFFFF1;
    // rom_array[34249] = 32'hFFFFFFF1;
    // rom_array[34250] = 32'hFFFFFFF1;
    // rom_array[34251] = 32'hFFFFFFF1;
    // rom_array[34252] = 32'hFFFFFFF1;
    // rom_array[34253] = 32'hFFFFFFF1;
    // rom_array[34254] = 32'hFFFFFFF1;
    // rom_array[34255] = 32'hFFFFFFF1;
    // rom_array[34256] = 32'hFFFFFFF1;
    // rom_array[34257] = 32'hFFFFFFF1;
    // rom_array[34258] = 32'hFFFFFFF1;
    // rom_array[34259] = 32'hFFFFFFF1;
    // rom_array[34260] = 32'hFFFFFFF1;
    // rom_array[34261] = 32'hFFFFFFF1;
    // rom_array[34262] = 32'hFFFFFFF1;
    // rom_array[34263] = 32'hFFFFFFF1;
    // rom_array[34264] = 32'hFFFFFFF1;
    // rom_array[34265] = 32'hFFFFFFF1;
    // rom_array[34266] = 32'hFFFFFFF1;
    // rom_array[34267] = 32'hFFFFFFF1;
    // rom_array[34268] = 32'hFFFFFFF1;
    // rom_array[34269] = 32'hFFFFFFF0;
    // rom_array[34270] = 32'hFFFFFFF0;
    // rom_array[34271] = 32'hFFFFFFF0;
    // rom_array[34272] = 32'hFFFFFFF0;
    // rom_array[34273] = 32'hFFFFFFF1;
    // rom_array[34274] = 32'hFFFFFFF1;
    // rom_array[34275] = 32'hFFFFFFF1;
    // rom_array[34276] = 32'hFFFFFFF1;
    // rom_array[34277] = 32'hFFFFFFF0;
    // rom_array[34278] = 32'hFFFFFFF0;
    // rom_array[34279] = 32'hFFFFFFF0;
    // rom_array[34280] = 32'hFFFFFFF0;
    // rom_array[34281] = 32'hFFFFFFF1;
    // rom_array[34282] = 32'hFFFFFFF1;
    // rom_array[34283] = 32'hFFFFFFF1;
    // rom_array[34284] = 32'hFFFFFFF1;
    // rom_array[34285] = 32'hFFFFFFF0;
    // rom_array[34286] = 32'hFFFFFFF0;
    // rom_array[34287] = 32'hFFFFFFF0;
    // rom_array[34288] = 32'hFFFFFFF0;
    // rom_array[34289] = 32'hFFFFFFF1;
    // rom_array[34290] = 32'hFFFFFFF1;
    // rom_array[34291] = 32'hFFFFFFF1;
    // rom_array[34292] = 32'hFFFFFFF1;
    // rom_array[34293] = 32'hFFFFFFF0;
    // rom_array[34294] = 32'hFFFFFFF0;
    // rom_array[34295] = 32'hFFFFFFF0;
    // rom_array[34296] = 32'hFFFFFFF0;
    // rom_array[34297] = 32'hFFFFFFF1;
    // rom_array[34298] = 32'hFFFFFFF1;
    // rom_array[34299] = 32'hFFFFFFF1;
    // rom_array[34300] = 32'hFFFFFFF1;
    // rom_array[34301] = 32'hFFFFFFF0;
    // rom_array[34302] = 32'hFFFFFFF0;
    // rom_array[34303] = 32'hFFFFFFF0;
    // rom_array[34304] = 32'hFFFFFFF0;
    // rom_array[34305] = 32'hFFFFFFF1;
    // rom_array[34306] = 32'hFFFFFFF1;
    // rom_array[34307] = 32'hFFFFFFF1;
    // rom_array[34308] = 32'hFFFFFFF1;
    // rom_array[34309] = 32'hFFFFFFF0;
    // rom_array[34310] = 32'hFFFFFFF0;
    // rom_array[34311] = 32'hFFFFFFF0;
    // rom_array[34312] = 32'hFFFFFFF0;
    // rom_array[34313] = 32'hFFFFFFF1;
    // rom_array[34314] = 32'hFFFFFFF1;
    // rom_array[34315] = 32'hFFFFFFF1;
    // rom_array[34316] = 32'hFFFFFFF1;
    // rom_array[34317] = 32'hFFFFFFF0;
    // rom_array[34318] = 32'hFFFFFFF0;
    // rom_array[34319] = 32'hFFFFFFF0;
    // rom_array[34320] = 32'hFFFFFFF0;
    // rom_array[34321] = 32'hFFFFFFF1;
    // rom_array[34322] = 32'hFFFFFFF1;
    // rom_array[34323] = 32'hFFFFFFF1;
    // rom_array[34324] = 32'hFFFFFFF1;
    // rom_array[34325] = 32'hFFFFFFF0;
    // rom_array[34326] = 32'hFFFFFFF0;
    // rom_array[34327] = 32'hFFFFFFF0;
    // rom_array[34328] = 32'hFFFFFFF0;
    // rom_array[34329] = 32'hFFFFFFF1;
    // rom_array[34330] = 32'hFFFFFFF1;
    // rom_array[34331] = 32'hFFFFFFF1;
    // rom_array[34332] = 32'hFFFFFFF1;
    // rom_array[34333] = 32'hFFFFFFF1;
    // rom_array[34334] = 32'hFFFFFFF1;
    // rom_array[34335] = 32'hFFFFFFF1;
    // rom_array[34336] = 32'hFFFFFFF1;
    // rom_array[34337] = 32'hFFFFFFF1;
    // rom_array[34338] = 32'hFFFFFFF1;
    // rom_array[34339] = 32'hFFFFFFF1;
    // rom_array[34340] = 32'hFFFFFFF1;
    // rom_array[34341] = 32'hFFFFFFF1;
    // rom_array[34342] = 32'hFFFFFFF1;
    // rom_array[34343] = 32'hFFFFFFF1;
    // rom_array[34344] = 32'hFFFFFFF1;
    // rom_array[34345] = 32'hFFFFFFF1;
    // rom_array[34346] = 32'hFFFFFFF1;
    // rom_array[34347] = 32'hFFFFFFF1;
    // rom_array[34348] = 32'hFFFFFFF1;
    // rom_array[34349] = 32'hFFFFFFF1;
    // rom_array[34350] = 32'hFFFFFFF1;
    // rom_array[34351] = 32'hFFFFFFF1;
    // rom_array[34352] = 32'hFFFFFFF1;
    // rom_array[34353] = 32'hFFFFFFF1;
    // rom_array[34354] = 32'hFFFFFFF1;
    // rom_array[34355] = 32'hFFFFFFF1;
    // rom_array[34356] = 32'hFFFFFFF1;
    // rom_array[34357] = 32'hFFFFFFF1;
    // rom_array[34358] = 32'hFFFFFFF1;
    // rom_array[34359] = 32'hFFFFFFF1;
    // rom_array[34360] = 32'hFFFFFFF1;
    // rom_array[34361] = 32'hFFFFFFF1;
    // rom_array[34362] = 32'hFFFFFFF1;
    // rom_array[34363] = 32'hFFFFFFF1;
    // rom_array[34364] = 32'hFFFFFFF1;
    // rom_array[34365] = 32'hFFFFFFF1;
    // rom_array[34366] = 32'hFFFFFFF1;
    // rom_array[34367] = 32'hFFFFFFF1;
    // rom_array[34368] = 32'hFFFFFFF1;
    // rom_array[34369] = 32'hFFFFFFF1;
    // rom_array[34370] = 32'hFFFFFFF1;
    // rom_array[34371] = 32'hFFFFFFF1;
    // rom_array[34372] = 32'hFFFFFFF1;
    // rom_array[34373] = 32'hFFFFFFF1;
    // rom_array[34374] = 32'hFFFFFFF1;
    // rom_array[34375] = 32'hFFFFFFF1;
    // rom_array[34376] = 32'hFFFFFFF1;
    // rom_array[34377] = 32'hFFFFFFF1;
    // rom_array[34378] = 32'hFFFFFFF1;
    // rom_array[34379] = 32'hFFFFFFF1;
    // rom_array[34380] = 32'hFFFFFFF1;
    // rom_array[34381] = 32'hFFFFFFF1;
    // rom_array[34382] = 32'hFFFFFFF1;
    // rom_array[34383] = 32'hFFFFFFF1;
    // rom_array[34384] = 32'hFFFFFFF1;
    // rom_array[34385] = 32'hFFFFFFF1;
    // rom_array[34386] = 32'hFFFFFFF1;
    // rom_array[34387] = 32'hFFFFFFF1;
    // rom_array[34388] = 32'hFFFFFFF1;
    // rom_array[34389] = 32'hFFFFFFF1;
    // rom_array[34390] = 32'hFFFFFFF1;
    // rom_array[34391] = 32'hFFFFFFF1;
    // rom_array[34392] = 32'hFFFFFFF1;
    // rom_array[34393] = 32'hFFFFFFF0;
    // rom_array[34394] = 32'hFFFFFFF0;
    // rom_array[34395] = 32'hFFFFFFF1;
    // rom_array[34396] = 32'hFFFFFFF1;
    // rom_array[34397] = 32'hFFFFFFF0;
    // rom_array[34398] = 32'hFFFFFFF0;
    // rom_array[34399] = 32'hFFFFFFF1;
    // rom_array[34400] = 32'hFFFFFFF1;
    // rom_array[34401] = 32'hFFFFFFF0;
    // rom_array[34402] = 32'hFFFFFFF0;
    // rom_array[34403] = 32'hFFFFFFF1;
    // rom_array[34404] = 32'hFFFFFFF1;
    // rom_array[34405] = 32'hFFFFFFF0;
    // rom_array[34406] = 32'hFFFFFFF0;
    // rom_array[34407] = 32'hFFFFFFF1;
    // rom_array[34408] = 32'hFFFFFFF1;
    // rom_array[34409] = 32'hFFFFFFF0;
    // rom_array[34410] = 32'hFFFFFFF0;
    // rom_array[34411] = 32'hFFFFFFF1;
    // rom_array[34412] = 32'hFFFFFFF1;
    // rom_array[34413] = 32'hFFFFFFF0;
    // rom_array[34414] = 32'hFFFFFFF0;
    // rom_array[34415] = 32'hFFFFFFF1;
    // rom_array[34416] = 32'hFFFFFFF1;
    // rom_array[34417] = 32'hFFFFFFF0;
    // rom_array[34418] = 32'hFFFFFFF0;
    // rom_array[34419] = 32'hFFFFFFF1;
    // rom_array[34420] = 32'hFFFFFFF1;
    // rom_array[34421] = 32'hFFFFFFF0;
    // rom_array[34422] = 32'hFFFFFFF0;
    // rom_array[34423] = 32'hFFFFFFF1;
    // rom_array[34424] = 32'hFFFFFFF1;
    // rom_array[34425] = 32'hFFFFFFF0;
    // rom_array[34426] = 32'hFFFFFFF0;
    // rom_array[34427] = 32'hFFFFFFF1;
    // rom_array[34428] = 32'hFFFFFFF1;
    // rom_array[34429] = 32'hFFFFFFF0;
    // rom_array[34430] = 32'hFFFFFFF0;
    // rom_array[34431] = 32'hFFFFFFF0;
    // rom_array[34432] = 32'hFFFFFFF0;
    // rom_array[34433] = 32'hFFFFFFF0;
    // rom_array[34434] = 32'hFFFFFFF0;
    // rom_array[34435] = 32'hFFFFFFF1;
    // rom_array[34436] = 32'hFFFFFFF1;
    // rom_array[34437] = 32'hFFFFFFF0;
    // rom_array[34438] = 32'hFFFFFFF0;
    // rom_array[34439] = 32'hFFFFFFF0;
    // rom_array[34440] = 32'hFFFFFFF0;
    // rom_array[34441] = 32'hFFFFFFF1;
    // rom_array[34442] = 32'hFFFFFFF1;
    // rom_array[34443] = 32'hFFFFFFF1;
    // rom_array[34444] = 32'hFFFFFFF1;
    // rom_array[34445] = 32'hFFFFFFF0;
    // rom_array[34446] = 32'hFFFFFFF0;
    // rom_array[34447] = 32'hFFFFFFF0;
    // rom_array[34448] = 32'hFFFFFFF0;
    // rom_array[34449] = 32'hFFFFFFF1;
    // rom_array[34450] = 32'hFFFFFFF1;
    // rom_array[34451] = 32'hFFFFFFF1;
    // rom_array[34452] = 32'hFFFFFFF1;
    // rom_array[34453] = 32'hFFFFFFF0;
    // rom_array[34454] = 32'hFFFFFFF0;
    // rom_array[34455] = 32'hFFFFFFF0;
    // rom_array[34456] = 32'hFFFFFFF0;
    // rom_array[34457] = 32'hFFFFFFF1;
    // rom_array[34458] = 32'hFFFFFFF1;
    // rom_array[34459] = 32'hFFFFFFF1;
    // rom_array[34460] = 32'hFFFFFFF1;
    // rom_array[34461] = 32'hFFFFFFF0;
    // rom_array[34462] = 32'hFFFFFFF0;
    // rom_array[34463] = 32'hFFFFFFF0;
    // rom_array[34464] = 32'hFFFFFFF0;
    // rom_array[34465] = 32'hFFFFFFF1;
    // rom_array[34466] = 32'hFFFFFFF1;
    // rom_array[34467] = 32'hFFFFFFF1;
    // rom_array[34468] = 32'hFFFFFFF1;
    // rom_array[34469] = 32'hFFFFFFF0;
    // rom_array[34470] = 32'hFFFFFFF0;
    // rom_array[34471] = 32'hFFFFFFF0;
    // rom_array[34472] = 32'hFFFFFFF0;
    // rom_array[34473] = 32'hFFFFFFF1;
    // rom_array[34474] = 32'hFFFFFFF1;
    // rom_array[34475] = 32'hFFFFFFF1;
    // rom_array[34476] = 32'hFFFFFFF1;
    // rom_array[34477] = 32'hFFFFFFF0;
    // rom_array[34478] = 32'hFFFFFFF0;
    // rom_array[34479] = 32'hFFFFFFF0;
    // rom_array[34480] = 32'hFFFFFFF0;
    // rom_array[34481] = 32'hFFFFFFF1;
    // rom_array[34482] = 32'hFFFFFFF1;
    // rom_array[34483] = 32'hFFFFFFF1;
    // rom_array[34484] = 32'hFFFFFFF1;
    // rom_array[34485] = 32'hFFFFFFF0;
    // rom_array[34486] = 32'hFFFFFFF0;
    // rom_array[34487] = 32'hFFFFFFF0;
    // rom_array[34488] = 32'hFFFFFFF0;
    // rom_array[34489] = 32'hFFFFFFF1;
    // rom_array[34490] = 32'hFFFFFFF1;
    // rom_array[34491] = 32'hFFFFFFF1;
    // rom_array[34492] = 32'hFFFFFFF1;
    // rom_array[34493] = 32'hFFFFFFF1;
    // rom_array[34494] = 32'hFFFFFFF1;
    // rom_array[34495] = 32'hFFFFFFF1;
    // rom_array[34496] = 32'hFFFFFFF1;
    // rom_array[34497] = 32'hFFFFFFF1;
    // rom_array[34498] = 32'hFFFFFFF1;
    // rom_array[34499] = 32'hFFFFFFF1;
    // rom_array[34500] = 32'hFFFFFFF1;
    // rom_array[34501] = 32'hFFFFFFF1;
    // rom_array[34502] = 32'hFFFFFFF1;
    // rom_array[34503] = 32'hFFFFFFF1;
    // rom_array[34504] = 32'hFFFFFFF1;
    // rom_array[34505] = 32'hFFFFFFF1;
    // rom_array[34506] = 32'hFFFFFFF1;
    // rom_array[34507] = 32'hFFFFFFF1;
    // rom_array[34508] = 32'hFFFFFFF1;
    // rom_array[34509] = 32'hFFFFFFF1;
    // rom_array[34510] = 32'hFFFFFFF1;
    // rom_array[34511] = 32'hFFFFFFF1;
    // rom_array[34512] = 32'hFFFFFFF1;
    // rom_array[34513] = 32'hFFFFFFF1;
    // rom_array[34514] = 32'hFFFFFFF1;
    // rom_array[34515] = 32'hFFFFFFF1;
    // rom_array[34516] = 32'hFFFFFFF1;
    // rom_array[34517] = 32'hFFFFFFF1;
    // rom_array[34518] = 32'hFFFFFFF1;
    // rom_array[34519] = 32'hFFFFFFF1;
    // rom_array[34520] = 32'hFFFFFFF1;
    // rom_array[34521] = 32'hFFFFFFF1;
    // rom_array[34522] = 32'hFFFFFFF1;
    // rom_array[34523] = 32'hFFFFFFF1;
    // rom_array[34524] = 32'hFFFFFFF1;
    // rom_array[34525] = 32'hFFFFFFF0;
    // rom_array[34526] = 32'hFFFFFFF0;
    // rom_array[34527] = 32'hFFFFFFF0;
    // rom_array[34528] = 32'hFFFFFFF0;
    // rom_array[34529] = 32'hFFFFFFF1;
    // rom_array[34530] = 32'hFFFFFFF1;
    // rom_array[34531] = 32'hFFFFFFF1;
    // rom_array[34532] = 32'hFFFFFFF1;
    // rom_array[34533] = 32'hFFFFFFF0;
    // rom_array[34534] = 32'hFFFFFFF0;
    // rom_array[34535] = 32'hFFFFFFF0;
    // rom_array[34536] = 32'hFFFFFFF0;
    // rom_array[34537] = 32'hFFFFFFF0;
    // rom_array[34538] = 32'hFFFFFFF0;
    // rom_array[34539] = 32'hFFFFFFF1;
    // rom_array[34540] = 32'hFFFFFFF1;
    // rom_array[34541] = 32'hFFFFFFF0;
    // rom_array[34542] = 32'hFFFFFFF0;
    // rom_array[34543] = 32'hFFFFFFF0;
    // rom_array[34544] = 32'hFFFFFFF0;
    // rom_array[34545] = 32'hFFFFFFF0;
    // rom_array[34546] = 32'hFFFFFFF0;
    // rom_array[34547] = 32'hFFFFFFF1;
    // rom_array[34548] = 32'hFFFFFFF1;
    // rom_array[34549] = 32'hFFFFFFF0;
    // rom_array[34550] = 32'hFFFFFFF0;
    // rom_array[34551] = 32'hFFFFFFF0;
    // rom_array[34552] = 32'hFFFFFFF0;
    // rom_array[34553] = 32'hFFFFFFF1;
    // rom_array[34554] = 32'hFFFFFFF1;
    // rom_array[34555] = 32'hFFFFFFF1;
    // rom_array[34556] = 32'hFFFFFFF1;
    // rom_array[34557] = 32'hFFFFFFF0;
    // rom_array[34558] = 32'hFFFFFFF0;
    // rom_array[34559] = 32'hFFFFFFF0;
    // rom_array[34560] = 32'hFFFFFFF0;
    // rom_array[34561] = 32'hFFFFFFF1;
    // rom_array[34562] = 32'hFFFFFFF1;
    // rom_array[34563] = 32'hFFFFFFF1;
    // rom_array[34564] = 32'hFFFFFFF1;
    // rom_array[34565] = 32'hFFFFFFF0;
    // rom_array[34566] = 32'hFFFFFFF0;
    // rom_array[34567] = 32'hFFFFFFF0;
    // rom_array[34568] = 32'hFFFFFFF0;
    // rom_array[34569] = 32'hFFFFFFF1;
    // rom_array[34570] = 32'hFFFFFFF1;
    // rom_array[34571] = 32'hFFFFFFF1;
    // rom_array[34572] = 32'hFFFFFFF1;
    // rom_array[34573] = 32'hFFFFFFF0;
    // rom_array[34574] = 32'hFFFFFFF0;
    // rom_array[34575] = 32'hFFFFFFF0;
    // rom_array[34576] = 32'hFFFFFFF0;
    // rom_array[34577] = 32'hFFFFFFF1;
    // rom_array[34578] = 32'hFFFFFFF1;
    // rom_array[34579] = 32'hFFFFFFF1;
    // rom_array[34580] = 32'hFFFFFFF1;
    // rom_array[34581] = 32'hFFFFFFF0;
    // rom_array[34582] = 32'hFFFFFFF0;
    // rom_array[34583] = 32'hFFFFFFF0;
    // rom_array[34584] = 32'hFFFFFFF0;
    // rom_array[34585] = 32'hFFFFFFF1;
    // rom_array[34586] = 32'hFFFFFFF1;
    // rom_array[34587] = 32'hFFFFFFF1;
    // rom_array[34588] = 32'hFFFFFFF1;
    // rom_array[34589] = 32'hFFFFFFF0;
    // rom_array[34590] = 32'hFFFFFFF0;
    // rom_array[34591] = 32'hFFFFFFF0;
    // rom_array[34592] = 32'hFFFFFFF0;
    // rom_array[34593] = 32'hFFFFFFF1;
    // rom_array[34594] = 32'hFFFFFFF1;
    // rom_array[34595] = 32'hFFFFFFF1;
    // rom_array[34596] = 32'hFFFFFFF1;
    // rom_array[34597] = 32'hFFFFFFF0;
    // rom_array[34598] = 32'hFFFFFFF0;
    // rom_array[34599] = 32'hFFFFFFF0;
    // rom_array[34600] = 32'hFFFFFFF0;
    // rom_array[34601] = 32'hFFFFFFF1;
    // rom_array[34602] = 32'hFFFFFFF1;
    // rom_array[34603] = 32'hFFFFFFF1;
    // rom_array[34604] = 32'hFFFFFFF1;
    // rom_array[34605] = 32'hFFFFFFF0;
    // rom_array[34606] = 32'hFFFFFFF0;
    // rom_array[34607] = 32'hFFFFFFF0;
    // rom_array[34608] = 32'hFFFFFFF0;
    // rom_array[34609] = 32'hFFFFFFF1;
    // rom_array[34610] = 32'hFFFFFFF1;
    // rom_array[34611] = 32'hFFFFFFF1;
    // rom_array[34612] = 32'hFFFFFFF1;
    // rom_array[34613] = 32'hFFFFFFF0;
    // rom_array[34614] = 32'hFFFFFFF0;
    // rom_array[34615] = 32'hFFFFFFF0;
    // rom_array[34616] = 32'hFFFFFFF0;
    // rom_array[34617] = 32'hFFFFFFF0;
    // rom_array[34618] = 32'hFFFFFFF0;
    // rom_array[34619] = 32'hFFFFFFF1;
    // rom_array[34620] = 32'hFFFFFFF1;
    // rom_array[34621] = 32'hFFFFFFF0;
    // rom_array[34622] = 32'hFFFFFFF0;
    // rom_array[34623] = 32'hFFFFFFF0;
    // rom_array[34624] = 32'hFFFFFFF0;
    // rom_array[34625] = 32'hFFFFFFF0;
    // rom_array[34626] = 32'hFFFFFFF0;
    // rom_array[34627] = 32'hFFFFFFF1;
    // rom_array[34628] = 32'hFFFFFFF1;
    // rom_array[34629] = 32'hFFFFFFF0;
    // rom_array[34630] = 32'hFFFFFFF0;
    // rom_array[34631] = 32'hFFFFFFF0;
    // rom_array[34632] = 32'hFFFFFFF0;
    // rom_array[34633] = 32'hFFFFFFF1;
    // rom_array[34634] = 32'hFFFFFFF1;
    // rom_array[34635] = 32'hFFFFFFF1;
    // rom_array[34636] = 32'hFFFFFFF1;
    // rom_array[34637] = 32'hFFFFFFF0;
    // rom_array[34638] = 32'hFFFFFFF0;
    // rom_array[34639] = 32'hFFFFFFF0;
    // rom_array[34640] = 32'hFFFFFFF0;
    // rom_array[34641] = 32'hFFFFFFF1;
    // rom_array[34642] = 32'hFFFFFFF1;
    // rom_array[34643] = 32'hFFFFFFF1;
    // rom_array[34644] = 32'hFFFFFFF1;
    // rom_array[34645] = 32'hFFFFFFF0;
    // rom_array[34646] = 32'hFFFFFFF0;
    // rom_array[34647] = 32'hFFFFFFF0;
    // rom_array[34648] = 32'hFFFFFFF0;
    // rom_array[34649] = 32'hFFFFFFF1;
    // rom_array[34650] = 32'hFFFFFFF1;
    // rom_array[34651] = 32'hFFFFFFF1;
    // rom_array[34652] = 32'hFFFFFFF1;
    // rom_array[34653] = 32'hFFFFFFF0;
    // rom_array[34654] = 32'hFFFFFFF0;
    // rom_array[34655] = 32'hFFFFFFF0;
    // rom_array[34656] = 32'hFFFFFFF0;
    // rom_array[34657] = 32'hFFFFFFF1;
    // rom_array[34658] = 32'hFFFFFFF1;
    // rom_array[34659] = 32'hFFFFFFF1;
    // rom_array[34660] = 32'hFFFFFFF1;
    // rom_array[34661] = 32'hFFFFFFF0;
    // rom_array[34662] = 32'hFFFFFFF0;
    // rom_array[34663] = 32'hFFFFFFF0;
    // rom_array[34664] = 32'hFFFFFFF0;
    // rom_array[34665] = 32'hFFFFFFF0;
    // rom_array[34666] = 32'hFFFFFFF0;
    // rom_array[34667] = 32'hFFFFFFF0;
    // rom_array[34668] = 32'hFFFFFFF0;
    // rom_array[34669] = 32'hFFFFFFF0;
    // rom_array[34670] = 32'hFFFFFFF0;
    // rom_array[34671] = 32'hFFFFFFF1;
    // rom_array[34672] = 32'hFFFFFFF1;
    // rom_array[34673] = 32'hFFFFFFF0;
    // rom_array[34674] = 32'hFFFFFFF0;
    // rom_array[34675] = 32'hFFFFFFF0;
    // rom_array[34676] = 32'hFFFFFFF0;
    // rom_array[34677] = 32'hFFFFFFF0;
    // rom_array[34678] = 32'hFFFFFFF0;
    // rom_array[34679] = 32'hFFFFFFF1;
    // rom_array[34680] = 32'hFFFFFFF1;
    // rom_array[34681] = 32'hFFFFFFF0;
    // rom_array[34682] = 32'hFFFFFFF0;
    // rom_array[34683] = 32'hFFFFFFF0;
    // rom_array[34684] = 32'hFFFFFFF0;
    // rom_array[34685] = 32'hFFFFFFF1;
    // rom_array[34686] = 32'hFFFFFFF1;
    // rom_array[34687] = 32'hFFFFFFF1;
    // rom_array[34688] = 32'hFFFFFFF1;
    // rom_array[34689] = 32'hFFFFFFF0;
    // rom_array[34690] = 32'hFFFFFFF0;
    // rom_array[34691] = 32'hFFFFFFF0;
    // rom_array[34692] = 32'hFFFFFFF0;
    // rom_array[34693] = 32'hFFFFFFF1;
    // rom_array[34694] = 32'hFFFFFFF1;
    // rom_array[34695] = 32'hFFFFFFF1;
    // rom_array[34696] = 32'hFFFFFFF1;
    // rom_array[34697] = 32'hFFFFFFF0;
    // rom_array[34698] = 32'hFFFFFFF0;
    // rom_array[34699] = 32'hFFFFFFF1;
    // rom_array[34700] = 32'hFFFFFFF1;
    // rom_array[34701] = 32'hFFFFFFF0;
    // rom_array[34702] = 32'hFFFFFFF0;
    // rom_array[34703] = 32'hFFFFFFF1;
    // rom_array[34704] = 32'hFFFFFFF1;
    // rom_array[34705] = 32'hFFFFFFF0;
    // rom_array[34706] = 32'hFFFFFFF0;
    // rom_array[34707] = 32'hFFFFFFF1;
    // rom_array[34708] = 32'hFFFFFFF1;
    // rom_array[34709] = 32'hFFFFFFF0;
    // rom_array[34710] = 32'hFFFFFFF0;
    // rom_array[34711] = 32'hFFFFFFF1;
    // rom_array[34712] = 32'hFFFFFFF1;
    // rom_array[34713] = 32'hFFFFFFF0;
    // rom_array[34714] = 32'hFFFFFFF0;
    // rom_array[34715] = 32'hFFFFFFF0;
    // rom_array[34716] = 32'hFFFFFFF0;
    // rom_array[34717] = 32'hFFFFFFF1;
    // rom_array[34718] = 32'hFFFFFFF1;
    // rom_array[34719] = 32'hFFFFFFF1;
    // rom_array[34720] = 32'hFFFFFFF1;
    // rom_array[34721] = 32'hFFFFFFF0;
    // rom_array[34722] = 32'hFFFFFFF0;
    // rom_array[34723] = 32'hFFFFFFF0;
    // rom_array[34724] = 32'hFFFFFFF0;
    // rom_array[34725] = 32'hFFFFFFF1;
    // rom_array[34726] = 32'hFFFFFFF1;
    // rom_array[34727] = 32'hFFFFFFF1;
    // rom_array[34728] = 32'hFFFFFFF1;
    // rom_array[34729] = 32'hFFFFFFF0;
    // rom_array[34730] = 32'hFFFFFFF0;
    // rom_array[34731] = 32'hFFFFFFF0;
    // rom_array[34732] = 32'hFFFFFFF0;
    // rom_array[34733] = 32'hFFFFFFF1;
    // rom_array[34734] = 32'hFFFFFFF1;
    // rom_array[34735] = 32'hFFFFFFF1;
    // rom_array[34736] = 32'hFFFFFFF1;
    // rom_array[34737] = 32'hFFFFFFF0;
    // rom_array[34738] = 32'hFFFFFFF0;
    // rom_array[34739] = 32'hFFFFFFF0;
    // rom_array[34740] = 32'hFFFFFFF0;
    // rom_array[34741] = 32'hFFFFFFF1;
    // rom_array[34742] = 32'hFFFFFFF1;
    // rom_array[34743] = 32'hFFFFFFF1;
    // rom_array[34744] = 32'hFFFFFFF1;
    // rom_array[34745] = 32'hFFFFFFF0;
    // rom_array[34746] = 32'hFFFFFFF0;
    // rom_array[34747] = 32'hFFFFFFF1;
    // rom_array[34748] = 32'hFFFFFFF1;
    // rom_array[34749] = 32'hFFFFFFF0;
    // rom_array[34750] = 32'hFFFFFFF0;
    // rom_array[34751] = 32'hFFFFFFF1;
    // rom_array[34752] = 32'hFFFFFFF1;
    // rom_array[34753] = 32'hFFFFFFF0;
    // rom_array[34754] = 32'hFFFFFFF0;
    // rom_array[34755] = 32'hFFFFFFF1;
    // rom_array[34756] = 32'hFFFFFFF1;
    // rom_array[34757] = 32'hFFFFFFF0;
    // rom_array[34758] = 32'hFFFFFFF0;
    // rom_array[34759] = 32'hFFFFFFF1;
    // rom_array[34760] = 32'hFFFFFFF1;
    // rom_array[34761] = 32'hFFFFFFF0;
    // rom_array[34762] = 32'hFFFFFFF0;
    // rom_array[34763] = 32'hFFFFFFF1;
    // rom_array[34764] = 32'hFFFFFFF1;
    // rom_array[34765] = 32'hFFFFFFF0;
    // rom_array[34766] = 32'hFFFFFFF0;
    // rom_array[34767] = 32'hFFFFFFF1;
    // rom_array[34768] = 32'hFFFFFFF1;
    // rom_array[34769] = 32'hFFFFFFF0;
    // rom_array[34770] = 32'hFFFFFFF0;
    // rom_array[34771] = 32'hFFFFFFF1;
    // rom_array[34772] = 32'hFFFFFFF1;
    // rom_array[34773] = 32'hFFFFFFF0;
    // rom_array[34774] = 32'hFFFFFFF0;
    // rom_array[34775] = 32'hFFFFFFF1;
    // rom_array[34776] = 32'hFFFFFFF1;
    // rom_array[34777] = 32'hFFFFFFF0;
    // rom_array[34778] = 32'hFFFFFFF0;
    // rom_array[34779] = 32'hFFFFFFF1;
    // rom_array[34780] = 32'hFFFFFFF1;
    // rom_array[34781] = 32'hFFFFFFF0;
    // rom_array[34782] = 32'hFFFFFFF0;
    // rom_array[34783] = 32'hFFFFFFF0;
    // rom_array[34784] = 32'hFFFFFFF0;
    // rom_array[34785] = 32'hFFFFFFF0;
    // rom_array[34786] = 32'hFFFFFFF0;
    // rom_array[34787] = 32'hFFFFFFF1;
    // rom_array[34788] = 32'hFFFFFFF1;
    // rom_array[34789] = 32'hFFFFFFF0;
    // rom_array[34790] = 32'hFFFFFFF0;
    // rom_array[34791] = 32'hFFFFFFF0;
    // rom_array[34792] = 32'hFFFFFFF0;
    // rom_array[34793] = 32'hFFFFFFF1;
    // rom_array[34794] = 32'hFFFFFFF1;
    // rom_array[34795] = 32'hFFFFFFF1;
    // rom_array[34796] = 32'hFFFFFFF1;
    // rom_array[34797] = 32'hFFFFFFF0;
    // rom_array[34798] = 32'hFFFFFFF0;
    // rom_array[34799] = 32'hFFFFFFF0;
    // rom_array[34800] = 32'hFFFFFFF0;
    // rom_array[34801] = 32'hFFFFFFF1;
    // rom_array[34802] = 32'hFFFFFFF1;
    // rom_array[34803] = 32'hFFFFFFF1;
    // rom_array[34804] = 32'hFFFFFFF1;
    // rom_array[34805] = 32'hFFFFFFF0;
    // rom_array[34806] = 32'hFFFFFFF0;
    // rom_array[34807] = 32'hFFFFFFF0;
    // rom_array[34808] = 32'hFFFFFFF0;
    // rom_array[34809] = 32'hFFFFFFF1;
    // rom_array[34810] = 32'hFFFFFFF1;
    // rom_array[34811] = 32'hFFFFFFF1;
    // rom_array[34812] = 32'hFFFFFFF1;
    // rom_array[34813] = 32'hFFFFFFF0;
    // rom_array[34814] = 32'hFFFFFFF0;
    // rom_array[34815] = 32'hFFFFFFF0;
    // rom_array[34816] = 32'hFFFFFFF0;
    // rom_array[34817] = 32'hFFFFFFF1;
    // rom_array[34818] = 32'hFFFFFFF1;
    // rom_array[34819] = 32'hFFFFFFF1;
    // rom_array[34820] = 32'hFFFFFFF1;
    // rom_array[34821] = 32'hFFFFFFF0;
    // rom_array[34822] = 32'hFFFFFFF0;
    // rom_array[34823] = 32'hFFFFFFF0;
    // rom_array[34824] = 32'hFFFFFFF0;
    // rom_array[34825] = 32'hFFFFFFF1;
    // rom_array[34826] = 32'hFFFFFFF1;
    // rom_array[34827] = 32'hFFFFFFF1;
    // rom_array[34828] = 32'hFFFFFFF1;
    // rom_array[34829] = 32'hFFFFFFF0;
    // rom_array[34830] = 32'hFFFFFFF0;
    // rom_array[34831] = 32'hFFFFFFF0;
    // rom_array[34832] = 32'hFFFFFFF0;
    // rom_array[34833] = 32'hFFFFFFF1;
    // rom_array[34834] = 32'hFFFFFFF1;
    // rom_array[34835] = 32'hFFFFFFF1;
    // rom_array[34836] = 32'hFFFFFFF1;
    // rom_array[34837] = 32'hFFFFFFF0;
    // rom_array[34838] = 32'hFFFFFFF0;
    // rom_array[34839] = 32'hFFFFFFF0;
    // rom_array[34840] = 32'hFFFFFFF0;
    // rom_array[34841] = 32'hFFFFFFF0;
    // rom_array[34842] = 32'hFFFFFFF0;
    // rom_array[34843] = 32'hFFFFFFF0;
    // rom_array[34844] = 32'hFFFFFFF0;
    // rom_array[34845] = 32'hFFFFFFF1;
    // rom_array[34846] = 32'hFFFFFFF1;
    // rom_array[34847] = 32'hFFFFFFF1;
    // rom_array[34848] = 32'hFFFFFFF1;
    // rom_array[34849] = 32'hFFFFFFF0;
    // rom_array[34850] = 32'hFFFFFFF0;
    // rom_array[34851] = 32'hFFFFFFF0;
    // rom_array[34852] = 32'hFFFFFFF0;
    // rom_array[34853] = 32'hFFFFFFF1;
    // rom_array[34854] = 32'hFFFFFFF1;
    // rom_array[34855] = 32'hFFFFFFF1;
    // rom_array[34856] = 32'hFFFFFFF1;
    // rom_array[34857] = 32'hFFFFFFF0;
    // rom_array[34858] = 32'hFFFFFFF0;
    // rom_array[34859] = 32'hFFFFFFF0;
    // rom_array[34860] = 32'hFFFFFFF0;
    // rom_array[34861] = 32'hFFFFFFF1;
    // rom_array[34862] = 32'hFFFFFFF1;
    // rom_array[34863] = 32'hFFFFFFF1;
    // rom_array[34864] = 32'hFFFFFFF1;
    // rom_array[34865] = 32'hFFFFFFF0;
    // rom_array[34866] = 32'hFFFFFFF0;
    // rom_array[34867] = 32'hFFFFFFF0;
    // rom_array[34868] = 32'hFFFFFFF0;
    // rom_array[34869] = 32'hFFFFFFF1;
    // rom_array[34870] = 32'hFFFFFFF1;
    // rom_array[34871] = 32'hFFFFFFF1;
    // rom_array[34872] = 32'hFFFFFFF1;
    // rom_array[34873] = 32'hFFFFFFF0;
    // rom_array[34874] = 32'hFFFFFFF0;
    // rom_array[34875] = 32'hFFFFFFF0;
    // rom_array[34876] = 32'hFFFFFFF0;
    // rom_array[34877] = 32'hFFFFFFF1;
    // rom_array[34878] = 32'hFFFFFFF1;
    // rom_array[34879] = 32'hFFFFFFF1;
    // rom_array[34880] = 32'hFFFFFFF1;
    // rom_array[34881] = 32'hFFFFFFF0;
    // rom_array[34882] = 32'hFFFFFFF0;
    // rom_array[34883] = 32'hFFFFFFF0;
    // rom_array[34884] = 32'hFFFFFFF0;
    // rom_array[34885] = 32'hFFFFFFF1;
    // rom_array[34886] = 32'hFFFFFFF1;
    // rom_array[34887] = 32'hFFFFFFF1;
    // rom_array[34888] = 32'hFFFFFFF1;
    // rom_array[34889] = 32'hFFFFFFF0;
    // rom_array[34890] = 32'hFFFFFFF0;
    // rom_array[34891] = 32'hFFFFFFF0;
    // rom_array[34892] = 32'hFFFFFFF0;
    // rom_array[34893] = 32'hFFFFFFF1;
    // rom_array[34894] = 32'hFFFFFFF1;
    // rom_array[34895] = 32'hFFFFFFF1;
    // rom_array[34896] = 32'hFFFFFFF1;
    // rom_array[34897] = 32'hFFFFFFF0;
    // rom_array[34898] = 32'hFFFFFFF0;
    // rom_array[34899] = 32'hFFFFFFF0;
    // rom_array[34900] = 32'hFFFFFFF0;
    // rom_array[34901] = 32'hFFFFFFF1;
    // rom_array[34902] = 32'hFFFFFFF1;
    // rom_array[34903] = 32'hFFFFFFF1;
    // rom_array[34904] = 32'hFFFFFFF1;
    // rom_array[34905] = 32'hFFFFFFF0;
    // rom_array[34906] = 32'hFFFFFFF0;
    // rom_array[34907] = 32'hFFFFFFF0;
    // rom_array[34908] = 32'hFFFFFFF0;
    // rom_array[34909] = 32'hFFFFFFF1;
    // rom_array[34910] = 32'hFFFFFFF1;
    // rom_array[34911] = 32'hFFFFFFF1;
    // rom_array[34912] = 32'hFFFFFFF1;
    // rom_array[34913] = 32'hFFFFFFF0;
    // rom_array[34914] = 32'hFFFFFFF0;
    // rom_array[34915] = 32'hFFFFFFF0;
    // rom_array[34916] = 32'hFFFFFFF0;
    // rom_array[34917] = 32'hFFFFFFF1;
    // rom_array[34918] = 32'hFFFFFFF1;
    // rom_array[34919] = 32'hFFFFFFF1;
    // rom_array[34920] = 32'hFFFFFFF1;
    // rom_array[34921] = 32'hFFFFFFF0;
    // rom_array[34922] = 32'hFFFFFFF0;
    // rom_array[34923] = 32'hFFFFFFF0;
    // rom_array[34924] = 32'hFFFFFFF0;
    // rom_array[34925] = 32'hFFFFFFF1;
    // rom_array[34926] = 32'hFFFFFFF1;
    // rom_array[34927] = 32'hFFFFFFF1;
    // rom_array[34928] = 32'hFFFFFFF1;
    // rom_array[34929] = 32'hFFFFFFF0;
    // rom_array[34930] = 32'hFFFFFFF0;
    // rom_array[34931] = 32'hFFFFFFF0;
    // rom_array[34932] = 32'hFFFFFFF0;
    // rom_array[34933] = 32'hFFFFFFF1;
    // rom_array[34934] = 32'hFFFFFFF1;
    // rom_array[34935] = 32'hFFFFFFF1;
    // rom_array[34936] = 32'hFFFFFFF1;
    // rom_array[34937] = 32'hFFFFFFF0;
    // rom_array[34938] = 32'hFFFFFFF0;
    // rom_array[34939] = 32'hFFFFFFF0;
    // rom_array[34940] = 32'hFFFFFFF0;
    // rom_array[34941] = 32'hFFFFFFF1;
    // rom_array[34942] = 32'hFFFFFFF1;
    // rom_array[34943] = 32'hFFFFFFF1;
    // rom_array[34944] = 32'hFFFFFFF1;
    // rom_array[34945] = 32'hFFFFFFF0;
    // rom_array[34946] = 32'hFFFFFFF0;
    // rom_array[34947] = 32'hFFFFFFF0;
    // rom_array[34948] = 32'hFFFFFFF0;
    // rom_array[34949] = 32'hFFFFFFF1;
    // rom_array[34950] = 32'hFFFFFFF1;
    // rom_array[34951] = 32'hFFFFFFF1;
    // rom_array[34952] = 32'hFFFFFFF1;
    // rom_array[34953] = 32'hFFFFFFF0;
    // rom_array[34954] = 32'hFFFFFFF0;
    // rom_array[34955] = 32'hFFFFFFF0;
    // rom_array[34956] = 32'hFFFFFFF0;
    // rom_array[34957] = 32'hFFFFFFF1;
    // rom_array[34958] = 32'hFFFFFFF1;
    // rom_array[34959] = 32'hFFFFFFF1;
    // rom_array[34960] = 32'hFFFFFFF1;
    // rom_array[34961] = 32'hFFFFFFF0;
    // rom_array[34962] = 32'hFFFFFFF0;
    // rom_array[34963] = 32'hFFFFFFF0;
    // rom_array[34964] = 32'hFFFFFFF0;
    // rom_array[34965] = 32'hFFFFFFF1;
    // rom_array[34966] = 32'hFFFFFFF1;
    // rom_array[34967] = 32'hFFFFFFF1;
    // rom_array[34968] = 32'hFFFFFFF1;
    // rom_array[34969] = 32'hFFFFFFF1;
    // rom_array[34970] = 32'hFFFFFFF1;
    // rom_array[34971] = 32'hFFFFFFF1;
    // rom_array[34972] = 32'hFFFFFFF1;
    // rom_array[34973] = 32'hFFFFFFF0;
    // rom_array[34974] = 32'hFFFFFFF0;
    // rom_array[34975] = 32'hFFFFFFF0;
    // rom_array[34976] = 32'hFFFFFFF0;
    // rom_array[34977] = 32'hFFFFFFF1;
    // rom_array[34978] = 32'hFFFFFFF1;
    // rom_array[34979] = 32'hFFFFFFF1;
    // rom_array[34980] = 32'hFFFFFFF1;
    // rom_array[34981] = 32'hFFFFFFF0;
    // rom_array[34982] = 32'hFFFFFFF0;
    // rom_array[34983] = 32'hFFFFFFF0;
    // rom_array[34984] = 32'hFFFFFFF0;
    // rom_array[34985] = 32'hFFFFFFF1;
    // rom_array[34986] = 32'hFFFFFFF1;
    // rom_array[34987] = 32'hFFFFFFF1;
    // rom_array[34988] = 32'hFFFFFFF1;
    // rom_array[34989] = 32'hFFFFFFF0;
    // rom_array[34990] = 32'hFFFFFFF0;
    // rom_array[34991] = 32'hFFFFFFF0;
    // rom_array[34992] = 32'hFFFFFFF0;
    // rom_array[34993] = 32'hFFFFFFF1;
    // rom_array[34994] = 32'hFFFFFFF1;
    // rom_array[34995] = 32'hFFFFFFF1;
    // rom_array[34996] = 32'hFFFFFFF1;
    // rom_array[34997] = 32'hFFFFFFF0;
    // rom_array[34998] = 32'hFFFFFFF0;
    // rom_array[34999] = 32'hFFFFFFF0;
    // rom_array[35000] = 32'hFFFFFFF0;
    // rom_array[35001] = 32'hFFFFFFF1;
    // rom_array[35002] = 32'hFFFFFFF1;
    // rom_array[35003] = 32'hFFFFFFF1;
    // rom_array[35004] = 32'hFFFFFFF1;
    // rom_array[35005] = 32'hFFFFFFF0;
    // rom_array[35006] = 32'hFFFFFFF0;
    // rom_array[35007] = 32'hFFFFFFF0;
    // rom_array[35008] = 32'hFFFFFFF0;
    // rom_array[35009] = 32'hFFFFFFF1;
    // rom_array[35010] = 32'hFFFFFFF1;
    // rom_array[35011] = 32'hFFFFFFF1;
    // rom_array[35012] = 32'hFFFFFFF1;
    // rom_array[35013] = 32'hFFFFFFF0;
    // rom_array[35014] = 32'hFFFFFFF0;
    // rom_array[35015] = 32'hFFFFFFF0;
    // rom_array[35016] = 32'hFFFFFFF0;
    // rom_array[35017] = 32'hFFFFFFF1;
    // rom_array[35018] = 32'hFFFFFFF1;
    // rom_array[35019] = 32'hFFFFFFF1;
    // rom_array[35020] = 32'hFFFFFFF1;
    // rom_array[35021] = 32'hFFFFFFF0;
    // rom_array[35022] = 32'hFFFFFFF0;
    // rom_array[35023] = 32'hFFFFFFF0;
    // rom_array[35024] = 32'hFFFFFFF0;
    // rom_array[35025] = 32'hFFFFFFF1;
    // rom_array[35026] = 32'hFFFFFFF1;
    // rom_array[35027] = 32'hFFFFFFF1;
    // rom_array[35028] = 32'hFFFFFFF1;
    // rom_array[35029] = 32'hFFFFFFF0;
    // rom_array[35030] = 32'hFFFFFFF0;
    // rom_array[35031] = 32'hFFFFFFF0;
    // rom_array[35032] = 32'hFFFFFFF0;
    // rom_array[35033] = 32'hFFFFFFF1;
    // rom_array[35034] = 32'hFFFFFFF1;
    // rom_array[35035] = 32'hFFFFFFF1;
    // rom_array[35036] = 32'hFFFFFFF1;
    // rom_array[35037] = 32'hFFFFFFF0;
    // rom_array[35038] = 32'hFFFFFFF0;
    // rom_array[35039] = 32'hFFFFFFF1;
    // rom_array[35040] = 32'hFFFFFFF1;
    // rom_array[35041] = 32'hFFFFFFF1;
    // rom_array[35042] = 32'hFFFFFFF1;
    // rom_array[35043] = 32'hFFFFFFF1;
    // rom_array[35044] = 32'hFFFFFFF1;
    // rom_array[35045] = 32'hFFFFFFF0;
    // rom_array[35046] = 32'hFFFFFFF0;
    // rom_array[35047] = 32'hFFFFFFF1;
    // rom_array[35048] = 32'hFFFFFFF1;
    // rom_array[35049] = 32'hFFFFFFF1;
    // rom_array[35050] = 32'hFFFFFFF1;
    // rom_array[35051] = 32'hFFFFFFF1;
    // rom_array[35052] = 32'hFFFFFFF1;
    // rom_array[35053] = 32'hFFFFFFF1;
    // rom_array[35054] = 32'hFFFFFFF1;
    // rom_array[35055] = 32'hFFFFFFF1;
    // rom_array[35056] = 32'hFFFFFFF1;
    // rom_array[35057] = 32'hFFFFFFF1;
    // rom_array[35058] = 32'hFFFFFFF1;
    // rom_array[35059] = 32'hFFFFFFF1;
    // rom_array[35060] = 32'hFFFFFFF1;
    // rom_array[35061] = 32'hFFFFFFF1;
    // rom_array[35062] = 32'hFFFFFFF1;
    // rom_array[35063] = 32'hFFFFFFF1;
    // rom_array[35064] = 32'hFFFFFFF1;
    // rom_array[35065] = 32'hFFFFFFF0;
    // rom_array[35066] = 32'hFFFFFFF0;
    // rom_array[35067] = 32'hFFFFFFF1;
    // rom_array[35068] = 32'hFFFFFFF1;
    // rom_array[35069] = 32'hFFFFFFF0;
    // rom_array[35070] = 32'hFFFFFFF0;
    // rom_array[35071] = 32'hFFFFFFF1;
    // rom_array[35072] = 32'hFFFFFFF1;
    // rom_array[35073] = 32'hFFFFFFF0;
    // rom_array[35074] = 32'hFFFFFFF0;
    // rom_array[35075] = 32'hFFFFFFF1;
    // rom_array[35076] = 32'hFFFFFFF1;
    // rom_array[35077] = 32'hFFFFFFF0;
    // rom_array[35078] = 32'hFFFFFFF0;
    // rom_array[35079] = 32'hFFFFFFF1;
    // rom_array[35080] = 32'hFFFFFFF1;
    // rom_array[35081] = 32'hFFFFFFF1;
    // rom_array[35082] = 32'hFFFFFFF1;
    // rom_array[35083] = 32'hFFFFFFF1;
    // rom_array[35084] = 32'hFFFFFFF1;
    // rom_array[35085] = 32'hFFFFFFF1;
    // rom_array[35086] = 32'hFFFFFFF1;
    // rom_array[35087] = 32'hFFFFFFF1;
    // rom_array[35088] = 32'hFFFFFFF1;
    // rom_array[35089] = 32'hFFFFFFF1;
    // rom_array[35090] = 32'hFFFFFFF1;
    // rom_array[35091] = 32'hFFFFFFF1;
    // rom_array[35092] = 32'hFFFFFFF1;
    // rom_array[35093] = 32'hFFFFFFF1;
    // rom_array[35094] = 32'hFFFFFFF1;
    // rom_array[35095] = 32'hFFFFFFF1;
    // rom_array[35096] = 32'hFFFFFFF1;
    // rom_array[35097] = 32'hFFFFFFF1;
    // rom_array[35098] = 32'hFFFFFFF1;
    // rom_array[35099] = 32'hFFFFFFF1;
    // rom_array[35100] = 32'hFFFFFFF1;
    // rom_array[35101] = 32'hFFFFFFF1;
    // rom_array[35102] = 32'hFFFFFFF1;
    // rom_array[35103] = 32'hFFFFFFF1;
    // rom_array[35104] = 32'hFFFFFFF1;
    // rom_array[35105] = 32'hFFFFFFF1;
    // rom_array[35106] = 32'hFFFFFFF1;
    // rom_array[35107] = 32'hFFFFFFF1;
    // rom_array[35108] = 32'hFFFFFFF1;
    // rom_array[35109] = 32'hFFFFFFF1;
    // rom_array[35110] = 32'hFFFFFFF1;
    // rom_array[35111] = 32'hFFFFFFF1;
    // rom_array[35112] = 32'hFFFFFFF1;
    // rom_array[35113] = 32'hFFFFFFF0;
    // rom_array[35114] = 32'hFFFFFFF0;
    // rom_array[35115] = 32'hFFFFFFF1;
    // rom_array[35116] = 32'hFFFFFFF1;
    // rom_array[35117] = 32'hFFFFFFF0;
    // rom_array[35118] = 32'hFFFFFFF0;
    // rom_array[35119] = 32'hFFFFFFF1;
    // rom_array[35120] = 32'hFFFFFFF1;
    // rom_array[35121] = 32'hFFFFFFF0;
    // rom_array[35122] = 32'hFFFFFFF0;
    // rom_array[35123] = 32'hFFFFFFF1;
    // rom_array[35124] = 32'hFFFFFFF1;
    // rom_array[35125] = 32'hFFFFFFF0;
    // rom_array[35126] = 32'hFFFFFFF0;
    // rom_array[35127] = 32'hFFFFFFF1;
    // rom_array[35128] = 32'hFFFFFFF1;
    // rom_array[35129] = 32'hFFFFFFF1;
    // rom_array[35130] = 32'hFFFFFFF1;
    // rom_array[35131] = 32'hFFFFFFF1;
    // rom_array[35132] = 32'hFFFFFFF1;
    // rom_array[35133] = 32'hFFFFFFF1;
    // rom_array[35134] = 32'hFFFFFFF1;
    // rom_array[35135] = 32'hFFFFFFF1;
    // rom_array[35136] = 32'hFFFFFFF1;
    // rom_array[35137] = 32'hFFFFFFF1;
    // rom_array[35138] = 32'hFFFFFFF1;
    // rom_array[35139] = 32'hFFFFFFF1;
    // rom_array[35140] = 32'hFFFFFFF1;
    // rom_array[35141] = 32'hFFFFFFF1;
    // rom_array[35142] = 32'hFFFFFFF1;
    // rom_array[35143] = 32'hFFFFFFF1;
    // rom_array[35144] = 32'hFFFFFFF1;
    // rom_array[35145] = 32'hFFFFFFF0;
    // rom_array[35146] = 32'hFFFFFFF0;
    // rom_array[35147] = 32'hFFFFFFF1;
    // rom_array[35148] = 32'hFFFFFFF1;
    // rom_array[35149] = 32'hFFFFFFF0;
    // rom_array[35150] = 32'hFFFFFFF0;
    // rom_array[35151] = 32'hFFFFFFF1;
    // rom_array[35152] = 32'hFFFFFFF1;
    // rom_array[35153] = 32'hFFFFFFF0;
    // rom_array[35154] = 32'hFFFFFFF0;
    // rom_array[35155] = 32'hFFFFFFF1;
    // rom_array[35156] = 32'hFFFFFFF1;
    // rom_array[35157] = 32'hFFFFFFF0;
    // rom_array[35158] = 32'hFFFFFFF0;
    // rom_array[35159] = 32'hFFFFFFF1;
    // rom_array[35160] = 32'hFFFFFFF1;
    // rom_array[35161] = 32'hFFFFFFF1;
    // rom_array[35162] = 32'hFFFFFFF1;
    // rom_array[35163] = 32'hFFFFFFF1;
    // rom_array[35164] = 32'hFFFFFFF1;
    // rom_array[35165] = 32'hFFFFFFF1;
    // rom_array[35166] = 32'hFFFFFFF1;
    // rom_array[35167] = 32'hFFFFFFF1;
    // rom_array[35168] = 32'hFFFFFFF1;
    // rom_array[35169] = 32'hFFFFFFF1;
    // rom_array[35170] = 32'hFFFFFFF1;
    // rom_array[35171] = 32'hFFFFFFF1;
    // rom_array[35172] = 32'hFFFFFFF1;
    // rom_array[35173] = 32'hFFFFFFF1;
    // rom_array[35174] = 32'hFFFFFFF1;
    // rom_array[35175] = 32'hFFFFFFF1;
    // rom_array[35176] = 32'hFFFFFFF1;
    // rom_array[35177] = 32'hFFFFFFF1;
    // rom_array[35178] = 32'hFFFFFFF1;
    // rom_array[35179] = 32'hFFFFFFF1;
    // rom_array[35180] = 32'hFFFFFFF1;
    // rom_array[35181] = 32'hFFFFFFF1;
    // rom_array[35182] = 32'hFFFFFFF1;
    // rom_array[35183] = 32'hFFFFFFF1;
    // rom_array[35184] = 32'hFFFFFFF1;
    // rom_array[35185] = 32'hFFFFFFF1;
    // rom_array[35186] = 32'hFFFFFFF1;
    // rom_array[35187] = 32'hFFFFFFF1;
    // rom_array[35188] = 32'hFFFFFFF1;
    // rom_array[35189] = 32'hFFFFFFF1;
    // rom_array[35190] = 32'hFFFFFFF1;
    // rom_array[35191] = 32'hFFFFFFF1;
    // rom_array[35192] = 32'hFFFFFFF1;
    // rom_array[35193] = 32'hFFFFFFF1;
    // rom_array[35194] = 32'hFFFFFFF1;
    // rom_array[35195] = 32'hFFFFFFF1;
    // rom_array[35196] = 32'hFFFFFFF1;
    // rom_array[35197] = 32'hFFFFFFF1;
    // rom_array[35198] = 32'hFFFFFFF1;
    // rom_array[35199] = 32'hFFFFFFF1;
    // rom_array[35200] = 32'hFFFFFFF1;
    // rom_array[35201] = 32'hFFFFFFF1;
    // rom_array[35202] = 32'hFFFFFFF1;
    // rom_array[35203] = 32'hFFFFFFF1;
    // rom_array[35204] = 32'hFFFFFFF1;
    // rom_array[35205] = 32'hFFFFFFF1;
    // rom_array[35206] = 32'hFFFFFFF1;
    // rom_array[35207] = 32'hFFFFFFF1;
    // rom_array[35208] = 32'hFFFFFFF1;
    // rom_array[35209] = 32'hFFFFFFF0;
    // rom_array[35210] = 32'hFFFFFFF0;
    // rom_array[35211] = 32'hFFFFFFF1;
    // rom_array[35212] = 32'hFFFFFFF1;
    // rom_array[35213] = 32'hFFFFFFF0;
    // rom_array[35214] = 32'hFFFFFFF0;
    // rom_array[35215] = 32'hFFFFFFF1;
    // rom_array[35216] = 32'hFFFFFFF1;
    // rom_array[35217] = 32'hFFFFFFF0;
    // rom_array[35218] = 32'hFFFFFFF0;
    // rom_array[35219] = 32'hFFFFFFF1;
    // rom_array[35220] = 32'hFFFFFFF1;
    // rom_array[35221] = 32'hFFFFFFF0;
    // rom_array[35222] = 32'hFFFFFFF0;
    // rom_array[35223] = 32'hFFFFFFF1;
    // rom_array[35224] = 32'hFFFFFFF1;
    // rom_array[35225] = 32'hFFFFFFF1;
    // rom_array[35226] = 32'hFFFFFFF1;
    // rom_array[35227] = 32'hFFFFFFF1;
    // rom_array[35228] = 32'hFFFFFFF1;
    // rom_array[35229] = 32'hFFFFFFF1;
    // rom_array[35230] = 32'hFFFFFFF1;
    // rom_array[35231] = 32'hFFFFFFF1;
    // rom_array[35232] = 32'hFFFFFFF1;
    // rom_array[35233] = 32'hFFFFFFF1;
    // rom_array[35234] = 32'hFFFFFFF1;
    // rom_array[35235] = 32'hFFFFFFF1;
    // rom_array[35236] = 32'hFFFFFFF1;
    // rom_array[35237] = 32'hFFFFFFF1;
    // rom_array[35238] = 32'hFFFFFFF1;
    // rom_array[35239] = 32'hFFFFFFF1;
    // rom_array[35240] = 32'hFFFFFFF1;
    // rom_array[35241] = 32'hFFFFFFF0;
    // rom_array[35242] = 32'hFFFFFFF0;
    // rom_array[35243] = 32'hFFFFFFF1;
    // rom_array[35244] = 32'hFFFFFFF1;
    // rom_array[35245] = 32'hFFFFFFF0;
    // rom_array[35246] = 32'hFFFFFFF0;
    // rom_array[35247] = 32'hFFFFFFF1;
    // rom_array[35248] = 32'hFFFFFFF1;
    // rom_array[35249] = 32'hFFFFFFF0;
    // rom_array[35250] = 32'hFFFFFFF0;
    // rom_array[35251] = 32'hFFFFFFF1;
    // rom_array[35252] = 32'hFFFFFFF1;
    // rom_array[35253] = 32'hFFFFFFF0;
    // rom_array[35254] = 32'hFFFFFFF0;
    // rom_array[35255] = 32'hFFFFFFF1;
    // rom_array[35256] = 32'hFFFFFFF1;
    // rom_array[35257] = 32'hFFFFFFF1;
    // rom_array[35258] = 32'hFFFFFFF1;
    // rom_array[35259] = 32'hFFFFFFF1;
    // rom_array[35260] = 32'hFFFFFFF1;
    // rom_array[35261] = 32'hFFFFFFF1;
    // rom_array[35262] = 32'hFFFFFFF1;
    // rom_array[35263] = 32'hFFFFFFF1;
    // rom_array[35264] = 32'hFFFFFFF1;
    // rom_array[35265] = 32'hFFFFFFF1;
    // rom_array[35266] = 32'hFFFFFFF1;
    // rom_array[35267] = 32'hFFFFFFF1;
    // rom_array[35268] = 32'hFFFFFFF1;
    // rom_array[35269] = 32'hFFFFFFF1;
    // rom_array[35270] = 32'hFFFFFFF1;
    // rom_array[35271] = 32'hFFFFFFF1;
    // rom_array[35272] = 32'hFFFFFFF1;
    // rom_array[35273] = 32'hFFFFFFF0;
    // rom_array[35274] = 32'hFFFFFFF0;
    // rom_array[35275] = 32'hFFFFFFF0;
    // rom_array[35276] = 32'hFFFFFFF0;
    // rom_array[35277] = 32'hFFFFFFF1;
    // rom_array[35278] = 32'hFFFFFFF1;
    // rom_array[35279] = 32'hFFFFFFF1;
    // rom_array[35280] = 32'hFFFFFFF1;
    // rom_array[35281] = 32'hFFFFFFF0;
    // rom_array[35282] = 32'hFFFFFFF0;
    // rom_array[35283] = 32'hFFFFFFF0;
    // rom_array[35284] = 32'hFFFFFFF0;
    // rom_array[35285] = 32'hFFFFFFF1;
    // rom_array[35286] = 32'hFFFFFFF1;
    // rom_array[35287] = 32'hFFFFFFF1;
    // rom_array[35288] = 32'hFFFFFFF1;
    // rom_array[35289] = 32'hFFFFFFF0;
    // rom_array[35290] = 32'hFFFFFFF0;
    // rom_array[35291] = 32'hFFFFFFF1;
    // rom_array[35292] = 32'hFFFFFFF1;
    // rom_array[35293] = 32'hFFFFFFF0;
    // rom_array[35294] = 32'hFFFFFFF0;
    // rom_array[35295] = 32'hFFFFFFF1;
    // rom_array[35296] = 32'hFFFFFFF1;
    // rom_array[35297] = 32'hFFFFFFF0;
    // rom_array[35298] = 32'hFFFFFFF0;
    // rom_array[35299] = 32'hFFFFFFF1;
    // rom_array[35300] = 32'hFFFFFFF1;
    // rom_array[35301] = 32'hFFFFFFF0;
    // rom_array[35302] = 32'hFFFFFFF0;
    // rom_array[35303] = 32'hFFFFFFF1;
    // rom_array[35304] = 32'hFFFFFFF1;
    // rom_array[35305] = 32'hFFFFFFF1;
    // rom_array[35306] = 32'hFFFFFFF1;
    // rom_array[35307] = 32'hFFFFFFF1;
    // rom_array[35308] = 32'hFFFFFFF1;
    // rom_array[35309] = 32'hFFFFFFF1;
    // rom_array[35310] = 32'hFFFFFFF1;
    // rom_array[35311] = 32'hFFFFFFF1;
    // rom_array[35312] = 32'hFFFFFFF1;
    // rom_array[35313] = 32'hFFFFFFF1;
    // rom_array[35314] = 32'hFFFFFFF1;
    // rom_array[35315] = 32'hFFFFFFF1;
    // rom_array[35316] = 32'hFFFFFFF1;
    // rom_array[35317] = 32'hFFFFFFF1;
    // rom_array[35318] = 32'hFFFFFFF1;
    // rom_array[35319] = 32'hFFFFFFF1;
    // rom_array[35320] = 32'hFFFFFFF1;
    // rom_array[35321] = 32'hFFFFFFF0;
    // rom_array[35322] = 32'hFFFFFFF0;
    // rom_array[35323] = 32'hFFFFFFF1;
    // rom_array[35324] = 32'hFFFFFFF1;
    // rom_array[35325] = 32'hFFFFFFF0;
    // rom_array[35326] = 32'hFFFFFFF0;
    // rom_array[35327] = 32'hFFFFFFF1;
    // rom_array[35328] = 32'hFFFFFFF1;
    // rom_array[35329] = 32'hFFFFFFF0;
    // rom_array[35330] = 32'hFFFFFFF0;
    // rom_array[35331] = 32'hFFFFFFF1;
    // rom_array[35332] = 32'hFFFFFFF1;
    // rom_array[35333] = 32'hFFFFFFF0;
    // rom_array[35334] = 32'hFFFFFFF0;
    // rom_array[35335] = 32'hFFFFFFF1;
    // rom_array[35336] = 32'hFFFFFFF1;
    // rom_array[35337] = 32'hFFFFFFF1;
    // rom_array[35338] = 32'hFFFFFFF1;
    // rom_array[35339] = 32'hFFFFFFF1;
    // rom_array[35340] = 32'hFFFFFFF1;
    // rom_array[35341] = 32'hFFFFFFF1;
    // rom_array[35342] = 32'hFFFFFFF1;
    // rom_array[35343] = 32'hFFFFFFF1;
    // rom_array[35344] = 32'hFFFFFFF1;
    // rom_array[35345] = 32'hFFFFFFF1;
    // rom_array[35346] = 32'hFFFFFFF1;
    // rom_array[35347] = 32'hFFFFFFF1;
    // rom_array[35348] = 32'hFFFFFFF1;
    // rom_array[35349] = 32'hFFFFFFF1;
    // rom_array[35350] = 32'hFFFFFFF1;
    // rom_array[35351] = 32'hFFFFFFF1;
    // rom_array[35352] = 32'hFFFFFFF1;
    // rom_array[35353] = 32'hFFFFFFF1;
    // rom_array[35354] = 32'hFFFFFFF1;
    // rom_array[35355] = 32'hFFFFFFF1;
    // rom_array[35356] = 32'hFFFFFFF1;
    // rom_array[35357] = 32'hFFFFFFF1;
    // rom_array[35358] = 32'hFFFFFFF1;
    // rom_array[35359] = 32'hFFFFFFF1;
    // rom_array[35360] = 32'hFFFFFFF1;
    // rom_array[35361] = 32'hFFFFFFF1;
    // rom_array[35362] = 32'hFFFFFFF1;
    // rom_array[35363] = 32'hFFFFFFF1;
    // rom_array[35364] = 32'hFFFFFFF1;
    // rom_array[35365] = 32'hFFFFFFF1;
    // rom_array[35366] = 32'hFFFFFFF1;
    // rom_array[35367] = 32'hFFFFFFF1;
    // rom_array[35368] = 32'hFFFFFFF1;
    // rom_array[35369] = 32'hFFFFFFF1;
    // rom_array[35370] = 32'hFFFFFFF1;
    // rom_array[35371] = 32'hFFFFFFF1;
    // rom_array[35372] = 32'hFFFFFFF1;
    // rom_array[35373] = 32'hFFFFFFF1;
    // rom_array[35374] = 32'hFFFFFFF1;
    // rom_array[35375] = 32'hFFFFFFF1;
    // rom_array[35376] = 32'hFFFFFFF1;
    // rom_array[35377] = 32'hFFFFFFF1;
    // rom_array[35378] = 32'hFFFFFFF1;
    // rom_array[35379] = 32'hFFFFFFF1;
    // rom_array[35380] = 32'hFFFFFFF1;
    // rom_array[35381] = 32'hFFFFFFF1;
    // rom_array[35382] = 32'hFFFFFFF1;
    // rom_array[35383] = 32'hFFFFFFF1;
    // rom_array[35384] = 32'hFFFFFFF1;
    // rom_array[35385] = 32'hFFFFFFF1;
    // rom_array[35386] = 32'hFFFFFFF1;
    // rom_array[35387] = 32'hFFFFFFF1;
    // rom_array[35388] = 32'hFFFFFFF1;
    // rom_array[35389] = 32'hFFFFFFF1;
    // rom_array[35390] = 32'hFFFFFFF1;
    // rom_array[35391] = 32'hFFFFFFF1;
    // rom_array[35392] = 32'hFFFFFFF1;
    // rom_array[35393] = 32'hFFFFFFF1;
    // rom_array[35394] = 32'hFFFFFFF1;
    // rom_array[35395] = 32'hFFFFFFF1;
    // rom_array[35396] = 32'hFFFFFFF1;
    // rom_array[35397] = 32'hFFFFFFF1;
    // rom_array[35398] = 32'hFFFFFFF1;
    // rom_array[35399] = 32'hFFFFFFF1;
    // rom_array[35400] = 32'hFFFFFFF1;
    // rom_array[35401] = 32'hFFFFFFF1;
    // rom_array[35402] = 32'hFFFFFFF1;
    // rom_array[35403] = 32'hFFFFFFF1;
    // rom_array[35404] = 32'hFFFFFFF1;
    // rom_array[35405] = 32'hFFFFFFF1;
    // rom_array[35406] = 32'hFFFFFFF1;
    // rom_array[35407] = 32'hFFFFFFF1;
    // rom_array[35408] = 32'hFFFFFFF1;
    // rom_array[35409] = 32'hFFFFFFF1;
    // rom_array[35410] = 32'hFFFFFFF1;
    // rom_array[35411] = 32'hFFFFFFF1;
    // rom_array[35412] = 32'hFFFFFFF1;
    // rom_array[35413] = 32'hFFFFFFF1;
    // rom_array[35414] = 32'hFFFFFFF1;
    // rom_array[35415] = 32'hFFFFFFF1;
    // rom_array[35416] = 32'hFFFFFFF1;
    // rom_array[35417] = 32'hFFFFFFF1;
    // rom_array[35418] = 32'hFFFFFFF1;
    // rom_array[35419] = 32'hFFFFFFF1;
    // rom_array[35420] = 32'hFFFFFFF1;
    // rom_array[35421] = 32'hFFFFFFF1;
    // rom_array[35422] = 32'hFFFFFFF1;
    // rom_array[35423] = 32'hFFFFFFF1;
    // rom_array[35424] = 32'hFFFFFFF1;
    // rom_array[35425] = 32'hFFFFFFF1;
    // rom_array[35426] = 32'hFFFFFFF1;
    // rom_array[35427] = 32'hFFFFFFF1;
    // rom_array[35428] = 32'hFFFFFFF1;
    // rom_array[35429] = 32'hFFFFFFF1;
    // rom_array[35430] = 32'hFFFFFFF1;
    // rom_array[35431] = 32'hFFFFFFF1;
    // rom_array[35432] = 32'hFFFFFFF1;
    // rom_array[35433] = 32'hFFFFFFF1;
    // rom_array[35434] = 32'hFFFFFFF1;
    // rom_array[35435] = 32'hFFFFFFF1;
    // rom_array[35436] = 32'hFFFFFFF1;
    // rom_array[35437] = 32'hFFFFFFF1;
    // rom_array[35438] = 32'hFFFFFFF1;
    // rom_array[35439] = 32'hFFFFFFF1;
    // rom_array[35440] = 32'hFFFFFFF1;
    // rom_array[35441] = 32'hFFFFFFF1;
    // rom_array[35442] = 32'hFFFFFFF1;
    // rom_array[35443] = 32'hFFFFFFF1;
    // rom_array[35444] = 32'hFFFFFFF1;
    // rom_array[35445] = 32'hFFFFFFF1;
    // rom_array[35446] = 32'hFFFFFFF1;
    // rom_array[35447] = 32'hFFFFFFF1;
    // rom_array[35448] = 32'hFFFFFFF1;
    // rom_array[35449] = 32'hFFFFFFF0;
    // rom_array[35450] = 32'hFFFFFFF0;
    // rom_array[35451] = 32'hFFFFFFF1;
    // rom_array[35452] = 32'hFFFFFFF1;
    // rom_array[35453] = 32'hFFFFFFF0;
    // rom_array[35454] = 32'hFFFFFFF0;
    // rom_array[35455] = 32'hFFFFFFF1;
    // rom_array[35456] = 32'hFFFFFFF1;
    // rom_array[35457] = 32'hFFFFFFF0;
    // rom_array[35458] = 32'hFFFFFFF0;
    // rom_array[35459] = 32'hFFFFFFF1;
    // rom_array[35460] = 32'hFFFFFFF1;
    // rom_array[35461] = 32'hFFFFFFF0;
    // rom_array[35462] = 32'hFFFFFFF0;
    // rom_array[35463] = 32'hFFFFFFF1;
    // rom_array[35464] = 32'hFFFFFFF1;
    // rom_array[35465] = 32'hFFFFFFF0;
    // rom_array[35466] = 32'hFFFFFFF0;
    // rom_array[35467] = 32'hFFFFFFF1;
    // rom_array[35468] = 32'hFFFFFFF1;
    // rom_array[35469] = 32'hFFFFFFF0;
    // rom_array[35470] = 32'hFFFFFFF0;
    // rom_array[35471] = 32'hFFFFFFF1;
    // rom_array[35472] = 32'hFFFFFFF1;
    // rom_array[35473] = 32'hFFFFFFF0;
    // rom_array[35474] = 32'hFFFFFFF0;
    // rom_array[35475] = 32'hFFFFFFF1;
    // rom_array[35476] = 32'hFFFFFFF1;
    // rom_array[35477] = 32'hFFFFFFF0;
    // rom_array[35478] = 32'hFFFFFFF0;
    // rom_array[35479] = 32'hFFFFFFF1;
    // rom_array[35480] = 32'hFFFFFFF1;
    // rom_array[35481] = 32'hFFFFFFF1;
    // rom_array[35482] = 32'hFFFFFFF1;
    // rom_array[35483] = 32'hFFFFFFF1;
    // rom_array[35484] = 32'hFFFFFFF1;
    // rom_array[35485] = 32'hFFFFFFF1;
    // rom_array[35486] = 32'hFFFFFFF1;
    // rom_array[35487] = 32'hFFFFFFF1;
    // rom_array[35488] = 32'hFFFFFFF1;
    // rom_array[35489] = 32'hFFFFFFF1;
    // rom_array[35490] = 32'hFFFFFFF1;
    // rom_array[35491] = 32'hFFFFFFF1;
    // rom_array[35492] = 32'hFFFFFFF1;
    // rom_array[35493] = 32'hFFFFFFF1;
    // rom_array[35494] = 32'hFFFFFFF1;
    // rom_array[35495] = 32'hFFFFFFF1;
    // rom_array[35496] = 32'hFFFFFFF1;
    // rom_array[35497] = 32'hFFFFFFF1;
    // rom_array[35498] = 32'hFFFFFFF1;
    // rom_array[35499] = 32'hFFFFFFF1;
    // rom_array[35500] = 32'hFFFFFFF1;
    // rom_array[35501] = 32'hFFFFFFF1;
    // rom_array[35502] = 32'hFFFFFFF1;
    // rom_array[35503] = 32'hFFFFFFF1;
    // rom_array[35504] = 32'hFFFFFFF1;
    // rom_array[35505] = 32'hFFFFFFF1;
    // rom_array[35506] = 32'hFFFFFFF1;
    // rom_array[35507] = 32'hFFFFFFF1;
    // rom_array[35508] = 32'hFFFFFFF1;
    // rom_array[35509] = 32'hFFFFFFF1;
    // rom_array[35510] = 32'hFFFFFFF1;
    // rom_array[35511] = 32'hFFFFFFF1;
    // rom_array[35512] = 32'hFFFFFFF1;
    // rom_array[35513] = 32'hFFFFFFF0;
    // rom_array[35514] = 32'hFFFFFFF0;
    // rom_array[35515] = 32'hFFFFFFF1;
    // rom_array[35516] = 32'hFFFFFFF1;
    // rom_array[35517] = 32'hFFFFFFF0;
    // rom_array[35518] = 32'hFFFFFFF0;
    // rom_array[35519] = 32'hFFFFFFF1;
    // rom_array[35520] = 32'hFFFFFFF1;
    // rom_array[35521] = 32'hFFFFFFF0;
    // rom_array[35522] = 32'hFFFFFFF0;
    // rom_array[35523] = 32'hFFFFFFF1;
    // rom_array[35524] = 32'hFFFFFFF1;
    // rom_array[35525] = 32'hFFFFFFF0;
    // rom_array[35526] = 32'hFFFFFFF0;
    // rom_array[35527] = 32'hFFFFFFF1;
    // rom_array[35528] = 32'hFFFFFFF1;
    // rom_array[35529] = 32'hFFFFFFF1;
    // rom_array[35530] = 32'hFFFFFFF1;
    // rom_array[35531] = 32'hFFFFFFF1;
    // rom_array[35532] = 32'hFFFFFFF1;
    // rom_array[35533] = 32'hFFFFFFF1;
    // rom_array[35534] = 32'hFFFFFFF1;
    // rom_array[35535] = 32'hFFFFFFF1;
    // rom_array[35536] = 32'hFFFFFFF1;
    // rom_array[35537] = 32'hFFFFFFF1;
    // rom_array[35538] = 32'hFFFFFFF1;
    // rom_array[35539] = 32'hFFFFFFF1;
    // rom_array[35540] = 32'hFFFFFFF1;
    // rom_array[35541] = 32'hFFFFFFF1;
    // rom_array[35542] = 32'hFFFFFFF1;
    // rom_array[35543] = 32'hFFFFFFF1;
    // rom_array[35544] = 32'hFFFFFFF1;
    // rom_array[35545] = 32'hFFFFFFF1;
    // rom_array[35546] = 32'hFFFFFFF1;
    // rom_array[35547] = 32'hFFFFFFF0;
    // rom_array[35548] = 32'hFFFFFFF0;
    // rom_array[35549] = 32'hFFFFFFF1;
    // rom_array[35550] = 32'hFFFFFFF1;
    // rom_array[35551] = 32'hFFFFFFF0;
    // rom_array[35552] = 32'hFFFFFFF0;
    // rom_array[35553] = 32'hFFFFFFF1;
    // rom_array[35554] = 32'hFFFFFFF1;
    // rom_array[35555] = 32'hFFFFFFF0;
    // rom_array[35556] = 32'hFFFFFFF0;
    // rom_array[35557] = 32'hFFFFFFF1;
    // rom_array[35558] = 32'hFFFFFFF1;
    // rom_array[35559] = 32'hFFFFFFF0;
    // rom_array[35560] = 32'hFFFFFFF0;
    // rom_array[35561] = 32'hFFFFFFF1;
    // rom_array[35562] = 32'hFFFFFFF1;
    // rom_array[35563] = 32'hFFFFFFF0;
    // rom_array[35564] = 32'hFFFFFFF0;
    // rom_array[35565] = 32'hFFFFFFF1;
    // rom_array[35566] = 32'hFFFFFFF1;
    // rom_array[35567] = 32'hFFFFFFF0;
    // rom_array[35568] = 32'hFFFFFFF0;
    // rom_array[35569] = 32'hFFFFFFF1;
    // rom_array[35570] = 32'hFFFFFFF1;
    // rom_array[35571] = 32'hFFFFFFF0;
    // rom_array[35572] = 32'hFFFFFFF0;
    // rom_array[35573] = 32'hFFFFFFF1;
    // rom_array[35574] = 32'hFFFFFFF1;
    // rom_array[35575] = 32'hFFFFFFF0;
    // rom_array[35576] = 32'hFFFFFFF0;
    // rom_array[35577] = 32'hFFFFFFF0;
    // rom_array[35578] = 32'hFFFFFFF0;
    // rom_array[35579] = 32'hFFFFFFF1;
    // rom_array[35580] = 32'hFFFFFFF1;
    // rom_array[35581] = 32'hFFFFFFF0;
    // rom_array[35582] = 32'hFFFFFFF0;
    // rom_array[35583] = 32'hFFFFFFF1;
    // rom_array[35584] = 32'hFFFFFFF1;
    // rom_array[35585] = 32'hFFFFFFF0;
    // rom_array[35586] = 32'hFFFFFFF0;
    // rom_array[35587] = 32'hFFFFFFF1;
    // rom_array[35588] = 32'hFFFFFFF1;
    // rom_array[35589] = 32'hFFFFFFF0;
    // rom_array[35590] = 32'hFFFFFFF0;
    // rom_array[35591] = 32'hFFFFFFF1;
    // rom_array[35592] = 32'hFFFFFFF1;
    // rom_array[35593] = 32'hFFFFFFF0;
    // rom_array[35594] = 32'hFFFFFFF0;
    // rom_array[35595] = 32'hFFFFFFF1;
    // rom_array[35596] = 32'hFFFFFFF1;
    // rom_array[35597] = 32'hFFFFFFF0;
    // rom_array[35598] = 32'hFFFFFFF0;
    // rom_array[35599] = 32'hFFFFFFF1;
    // rom_array[35600] = 32'hFFFFFFF1;
    // rom_array[35601] = 32'hFFFFFFF0;
    // rom_array[35602] = 32'hFFFFFFF0;
    // rom_array[35603] = 32'hFFFFFFF1;
    // rom_array[35604] = 32'hFFFFFFF1;
    // rom_array[35605] = 32'hFFFFFFF0;
    // rom_array[35606] = 32'hFFFFFFF0;
    // rom_array[35607] = 32'hFFFFFFF1;
    // rom_array[35608] = 32'hFFFFFFF1;
    // rom_array[35609] = 32'hFFFFFFF1;
    // rom_array[35610] = 32'hFFFFFFF1;
    // rom_array[35611] = 32'hFFFFFFF0;
    // rom_array[35612] = 32'hFFFFFFF0;
    // rom_array[35613] = 32'hFFFFFFF1;
    // rom_array[35614] = 32'hFFFFFFF1;
    // rom_array[35615] = 32'hFFFFFFF0;
    // rom_array[35616] = 32'hFFFFFFF0;
    // rom_array[35617] = 32'hFFFFFFF1;
    // rom_array[35618] = 32'hFFFFFFF1;
    // rom_array[35619] = 32'hFFFFFFF0;
    // rom_array[35620] = 32'hFFFFFFF0;
    // rom_array[35621] = 32'hFFFFFFF1;
    // rom_array[35622] = 32'hFFFFFFF1;
    // rom_array[35623] = 32'hFFFFFFF0;
    // rom_array[35624] = 32'hFFFFFFF0;
    // rom_array[35625] = 32'hFFFFFFF1;
    // rom_array[35626] = 32'hFFFFFFF1;
    // rom_array[35627] = 32'hFFFFFFF0;
    // rom_array[35628] = 32'hFFFFFFF0;
    // rom_array[35629] = 32'hFFFFFFF1;
    // rom_array[35630] = 32'hFFFFFFF1;
    // rom_array[35631] = 32'hFFFFFFF1;
    // rom_array[35632] = 32'hFFFFFFF1;
    // rom_array[35633] = 32'hFFFFFFF1;
    // rom_array[35634] = 32'hFFFFFFF1;
    // rom_array[35635] = 32'hFFFFFFF0;
    // rom_array[35636] = 32'hFFFFFFF0;
    // rom_array[35637] = 32'hFFFFFFF1;
    // rom_array[35638] = 32'hFFFFFFF1;
    // rom_array[35639] = 32'hFFFFFFF1;
    // rom_array[35640] = 32'hFFFFFFF1;
    // rom_array[35641] = 32'hFFFFFFF0;
    // rom_array[35642] = 32'hFFFFFFF0;
    // rom_array[35643] = 32'hFFFFFFF1;
    // rom_array[35644] = 32'hFFFFFFF1;
    // rom_array[35645] = 32'hFFFFFFF0;
    // rom_array[35646] = 32'hFFFFFFF0;
    // rom_array[35647] = 32'hFFFFFFF0;
    // rom_array[35648] = 32'hFFFFFFF0;
    // rom_array[35649] = 32'hFFFFFFF0;
    // rom_array[35650] = 32'hFFFFFFF0;
    // rom_array[35651] = 32'hFFFFFFF1;
    // rom_array[35652] = 32'hFFFFFFF1;
    // rom_array[35653] = 32'hFFFFFFF0;
    // rom_array[35654] = 32'hFFFFFFF0;
    // rom_array[35655] = 32'hFFFFFFF0;
    // rom_array[35656] = 32'hFFFFFFF0;
    // rom_array[35657] = 32'hFFFFFFF1;
    // rom_array[35658] = 32'hFFFFFFF1;
    // rom_array[35659] = 32'hFFFFFFF1;
    // rom_array[35660] = 32'hFFFFFFF1;
    // rom_array[35661] = 32'hFFFFFFF0;
    // rom_array[35662] = 32'hFFFFFFF0;
    // rom_array[35663] = 32'hFFFFFFF0;
    // rom_array[35664] = 32'hFFFFFFF0;
    // rom_array[35665] = 32'hFFFFFFF1;
    // rom_array[35666] = 32'hFFFFFFF1;
    // rom_array[35667] = 32'hFFFFFFF1;
    // rom_array[35668] = 32'hFFFFFFF1;
    // rom_array[35669] = 32'hFFFFFFF0;
    // rom_array[35670] = 32'hFFFFFFF0;
    // rom_array[35671] = 32'hFFFFFFF0;
    // rom_array[35672] = 32'hFFFFFFF0;
    // rom_array[35673] = 32'hFFFFFFF1;
    // rom_array[35674] = 32'hFFFFFFF1;
    // rom_array[35675] = 32'hFFFFFFF1;
    // rom_array[35676] = 32'hFFFFFFF1;
    // rom_array[35677] = 32'hFFFFFFF0;
    // rom_array[35678] = 32'hFFFFFFF0;
    // rom_array[35679] = 32'hFFFFFFF0;
    // rom_array[35680] = 32'hFFFFFFF0;
    // rom_array[35681] = 32'hFFFFFFF1;
    // rom_array[35682] = 32'hFFFFFFF1;
    // rom_array[35683] = 32'hFFFFFFF1;
    // rom_array[35684] = 32'hFFFFFFF1;
    // rom_array[35685] = 32'hFFFFFFF0;
    // rom_array[35686] = 32'hFFFFFFF0;
    // rom_array[35687] = 32'hFFFFFFF0;
    // rom_array[35688] = 32'hFFFFFFF0;
    // rom_array[35689] = 32'hFFFFFFF1;
    // rom_array[35690] = 32'hFFFFFFF1;
    // rom_array[35691] = 32'hFFFFFFF1;
    // rom_array[35692] = 32'hFFFFFFF1;
    // rom_array[35693] = 32'hFFFFFFF1;
    // rom_array[35694] = 32'hFFFFFFF1;
    // rom_array[35695] = 32'hFFFFFFF1;
    // rom_array[35696] = 32'hFFFFFFF1;
    // rom_array[35697] = 32'hFFFFFFF1;
    // rom_array[35698] = 32'hFFFFFFF1;
    // rom_array[35699] = 32'hFFFFFFF1;
    // rom_array[35700] = 32'hFFFFFFF1;
    // rom_array[35701] = 32'hFFFFFFF1;
    // rom_array[35702] = 32'hFFFFFFF1;
    // rom_array[35703] = 32'hFFFFFFF1;
    // rom_array[35704] = 32'hFFFFFFF1;
    // rom_array[35705] = 32'hFFFFFFF1;
    // rom_array[35706] = 32'hFFFFFFF1;
    // rom_array[35707] = 32'hFFFFFFF1;
    // rom_array[35708] = 32'hFFFFFFF1;
    // rom_array[35709] = 32'hFFFFFFF1;
    // rom_array[35710] = 32'hFFFFFFF1;
    // rom_array[35711] = 32'hFFFFFFF1;
    // rom_array[35712] = 32'hFFFFFFF1;
    // rom_array[35713] = 32'hFFFFFFF1;
    // rom_array[35714] = 32'hFFFFFFF1;
    // rom_array[35715] = 32'hFFFFFFF1;
    // rom_array[35716] = 32'hFFFFFFF1;
    // rom_array[35717] = 32'hFFFFFFF1;
    // rom_array[35718] = 32'hFFFFFFF1;
    // rom_array[35719] = 32'hFFFFFFF1;
    // rom_array[35720] = 32'hFFFFFFF1;
    // rom_array[35721] = 32'hFFFFFFF0;
    // rom_array[35722] = 32'hFFFFFFF0;
    // rom_array[35723] = 32'hFFFFFFF1;
    // rom_array[35724] = 32'hFFFFFFF1;
    // rom_array[35725] = 32'hFFFFFFF0;
    // rom_array[35726] = 32'hFFFFFFF0;
    // rom_array[35727] = 32'hFFFFFFF1;
    // rom_array[35728] = 32'hFFFFFFF1;
    // rom_array[35729] = 32'hFFFFFFF0;
    // rom_array[35730] = 32'hFFFFFFF0;
    // rom_array[35731] = 32'hFFFFFFF1;
    // rom_array[35732] = 32'hFFFFFFF1;
    // rom_array[35733] = 32'hFFFFFFF0;
    // rom_array[35734] = 32'hFFFFFFF0;
    // rom_array[35735] = 32'hFFFFFFF1;
    // rom_array[35736] = 32'hFFFFFFF1;
    // rom_array[35737] = 32'hFFFFFFF1;
    // rom_array[35738] = 32'hFFFFFFF1;
    // rom_array[35739] = 32'hFFFFFFF1;
    // rom_array[35740] = 32'hFFFFFFF1;
    // rom_array[35741] = 32'hFFFFFFF1;
    // rom_array[35742] = 32'hFFFFFFF1;
    // rom_array[35743] = 32'hFFFFFFF1;
    // rom_array[35744] = 32'hFFFFFFF1;
    // rom_array[35745] = 32'hFFFFFFF1;
    // rom_array[35746] = 32'hFFFFFFF1;
    // rom_array[35747] = 32'hFFFFFFF1;
    // rom_array[35748] = 32'hFFFFFFF1;
    // rom_array[35749] = 32'hFFFFFFF1;
    // rom_array[35750] = 32'hFFFFFFF1;
    // rom_array[35751] = 32'hFFFFFFF1;
    // rom_array[35752] = 32'hFFFFFFF1;
    // rom_array[35753] = 32'hFFFFFFF0;
    // rom_array[35754] = 32'hFFFFFFF0;
    // rom_array[35755] = 32'hFFFFFFF1;
    // rom_array[35756] = 32'hFFFFFFF1;
    // rom_array[35757] = 32'hFFFFFFF0;
    // rom_array[35758] = 32'hFFFFFFF0;
    // rom_array[35759] = 32'hFFFFFFF0;
    // rom_array[35760] = 32'hFFFFFFF0;
    // rom_array[35761] = 32'hFFFFFFF0;
    // rom_array[35762] = 32'hFFFFFFF0;
    // rom_array[35763] = 32'hFFFFFFF1;
    // rom_array[35764] = 32'hFFFFFFF1;
    // rom_array[35765] = 32'hFFFFFFF0;
    // rom_array[35766] = 32'hFFFFFFF0;
    // rom_array[35767] = 32'hFFFFFFF0;
    // rom_array[35768] = 32'hFFFFFFF0;
    // rom_array[35769] = 32'hFFFFFFF1;
    // rom_array[35770] = 32'hFFFFFFF1;
    // rom_array[35771] = 32'hFFFFFFF1;
    // rom_array[35772] = 32'hFFFFFFF1;
    // rom_array[35773] = 32'hFFFFFFF0;
    // rom_array[35774] = 32'hFFFFFFF0;
    // rom_array[35775] = 32'hFFFFFFF0;
    // rom_array[35776] = 32'hFFFFFFF0;
    // rom_array[35777] = 32'hFFFFFFF1;
    // rom_array[35778] = 32'hFFFFFFF1;
    // rom_array[35779] = 32'hFFFFFFF1;
    // rom_array[35780] = 32'hFFFFFFF1;
    // rom_array[35781] = 32'hFFFFFFF0;
    // rom_array[35782] = 32'hFFFFFFF0;
    // rom_array[35783] = 32'hFFFFFFF0;
    // rom_array[35784] = 32'hFFFFFFF0;
    // rom_array[35785] = 32'hFFFFFFF1;
    // rom_array[35786] = 32'hFFFFFFF1;
    // rom_array[35787] = 32'hFFFFFFF1;
    // rom_array[35788] = 32'hFFFFFFF1;
    // rom_array[35789] = 32'hFFFFFFF1;
    // rom_array[35790] = 32'hFFFFFFF1;
    // rom_array[35791] = 32'hFFFFFFF1;
    // rom_array[35792] = 32'hFFFFFFF1;
    // rom_array[35793] = 32'hFFFFFFF1;
    // rom_array[35794] = 32'hFFFFFFF1;
    // rom_array[35795] = 32'hFFFFFFF1;
    // rom_array[35796] = 32'hFFFFFFF1;
    // rom_array[35797] = 32'hFFFFFFF1;
    // rom_array[35798] = 32'hFFFFFFF1;
    // rom_array[35799] = 32'hFFFFFFF1;
    // rom_array[35800] = 32'hFFFFFFF1;
    // rom_array[35801] = 32'hFFFFFFF1;
    // rom_array[35802] = 32'hFFFFFFF1;
    // rom_array[35803] = 32'hFFFFFFF1;
    // rom_array[35804] = 32'hFFFFFFF1;
    // rom_array[35805] = 32'hFFFFFFF0;
    // rom_array[35806] = 32'hFFFFFFF0;
    // rom_array[35807] = 32'hFFFFFFF0;
    // rom_array[35808] = 32'hFFFFFFF0;
    // rom_array[35809] = 32'hFFFFFFF1;
    // rom_array[35810] = 32'hFFFFFFF1;
    // rom_array[35811] = 32'hFFFFFFF1;
    // rom_array[35812] = 32'hFFFFFFF1;
    // rom_array[35813] = 32'hFFFFFFF0;
    // rom_array[35814] = 32'hFFFFFFF0;
    // rom_array[35815] = 32'hFFFFFFF0;
    // rom_array[35816] = 32'hFFFFFFF0;
    // rom_array[35817] = 32'hFFFFFFF1;
    // rom_array[35818] = 32'hFFFFFFF1;
    // rom_array[35819] = 32'hFFFFFFF1;
    // rom_array[35820] = 32'hFFFFFFF1;
    // rom_array[35821] = 32'hFFFFFFF0;
    // rom_array[35822] = 32'hFFFFFFF0;
    // rom_array[35823] = 32'hFFFFFFF0;
    // rom_array[35824] = 32'hFFFFFFF0;
    // rom_array[35825] = 32'hFFFFFFF1;
    // rom_array[35826] = 32'hFFFFFFF1;
    // rom_array[35827] = 32'hFFFFFFF1;
    // rom_array[35828] = 32'hFFFFFFF1;
    // rom_array[35829] = 32'hFFFFFFF0;
    // rom_array[35830] = 32'hFFFFFFF0;
    // rom_array[35831] = 32'hFFFFFFF0;
    // rom_array[35832] = 32'hFFFFFFF0;
    // rom_array[35833] = 32'hFFFFFFF1;
    // rom_array[35834] = 32'hFFFFFFF1;
    // rom_array[35835] = 32'hFFFFFFF1;
    // rom_array[35836] = 32'hFFFFFFF1;
    // rom_array[35837] = 32'hFFFFFFF0;
    // rom_array[35838] = 32'hFFFFFFF0;
    // rom_array[35839] = 32'hFFFFFFF0;
    // rom_array[35840] = 32'hFFFFFFF0;
    // rom_array[35841] = 32'hFFFFFFF1;
    // rom_array[35842] = 32'hFFFFFFF1;
    // rom_array[35843] = 32'hFFFFFFF1;
    // rom_array[35844] = 32'hFFFFFFF1;
    // rom_array[35845] = 32'hFFFFFFF0;
    // rom_array[35846] = 32'hFFFFFFF0;
    // rom_array[35847] = 32'hFFFFFFF0;
    // rom_array[35848] = 32'hFFFFFFF0;
    // rom_array[35849] = 32'hFFFFFFF1;
    // rom_array[35850] = 32'hFFFFFFF1;
    // rom_array[35851] = 32'hFFFFFFF1;
    // rom_array[35852] = 32'hFFFFFFF1;
    // rom_array[35853] = 32'hFFFFFFF0;
    // rom_array[35854] = 32'hFFFFFFF0;
    // rom_array[35855] = 32'hFFFFFFF0;
    // rom_array[35856] = 32'hFFFFFFF0;
    // rom_array[35857] = 32'hFFFFFFF1;
    // rom_array[35858] = 32'hFFFFFFF1;
    // rom_array[35859] = 32'hFFFFFFF1;
    // rom_array[35860] = 32'hFFFFFFF1;
    // rom_array[35861] = 32'hFFFFFFF0;
    // rom_array[35862] = 32'hFFFFFFF0;
    // rom_array[35863] = 32'hFFFFFFF0;
    // rom_array[35864] = 32'hFFFFFFF0;
    // rom_array[35865] = 32'hFFFFFFF1;
    // rom_array[35866] = 32'hFFFFFFF1;
    // rom_array[35867] = 32'hFFFFFFF1;
    // rom_array[35868] = 32'hFFFFFFF1;
    // rom_array[35869] = 32'hFFFFFFF0;
    // rom_array[35870] = 32'hFFFFFFF0;
    // rom_array[35871] = 32'hFFFFFFF0;
    // rom_array[35872] = 32'hFFFFFFF0;
    // rom_array[35873] = 32'hFFFFFFF1;
    // rom_array[35874] = 32'hFFFFFFF1;
    // rom_array[35875] = 32'hFFFFFFF1;
    // rom_array[35876] = 32'hFFFFFFF1;
    // rom_array[35877] = 32'hFFFFFFF0;
    // rom_array[35878] = 32'hFFFFFFF0;
    // rom_array[35879] = 32'hFFFFFFF0;
    // rom_array[35880] = 32'hFFFFFFF0;
    // rom_array[35881] = 32'hFFFFFFF1;
    // rom_array[35882] = 32'hFFFFFFF1;
    // rom_array[35883] = 32'hFFFFFFF1;
    // rom_array[35884] = 32'hFFFFFFF1;
    // rom_array[35885] = 32'hFFFFFFF0;
    // rom_array[35886] = 32'hFFFFFFF0;
    // rom_array[35887] = 32'hFFFFFFF0;
    // rom_array[35888] = 32'hFFFFFFF0;
    // rom_array[35889] = 32'hFFFFFFF1;
    // rom_array[35890] = 32'hFFFFFFF1;
    // rom_array[35891] = 32'hFFFFFFF1;
    // rom_array[35892] = 32'hFFFFFFF1;
    // rom_array[35893] = 32'hFFFFFFF0;
    // rom_array[35894] = 32'hFFFFFFF0;
    // rom_array[35895] = 32'hFFFFFFF0;
    // rom_array[35896] = 32'hFFFFFFF0;
    // rom_array[35897] = 32'hFFFFFFF1;
    // rom_array[35898] = 32'hFFFFFFF1;
    // rom_array[35899] = 32'hFFFFFFF1;
    // rom_array[35900] = 32'hFFFFFFF1;
    // rom_array[35901] = 32'hFFFFFFF0;
    // rom_array[35902] = 32'hFFFFFFF0;
    // rom_array[35903] = 32'hFFFFFFF0;
    // rom_array[35904] = 32'hFFFFFFF0;
    // rom_array[35905] = 32'hFFFFFFF1;
    // rom_array[35906] = 32'hFFFFFFF1;
    // rom_array[35907] = 32'hFFFFFFF1;
    // rom_array[35908] = 32'hFFFFFFF1;
    // rom_array[35909] = 32'hFFFFFFF0;
    // rom_array[35910] = 32'hFFFFFFF0;
    // rom_array[35911] = 32'hFFFFFFF0;
    // rom_array[35912] = 32'hFFFFFFF0;
    // rom_array[35913] = 32'hFFFFFFF1;
    // rom_array[35914] = 32'hFFFFFFF1;
    // rom_array[35915] = 32'hFFFFFFF1;
    // rom_array[35916] = 32'hFFFFFFF1;
    // rom_array[35917] = 32'hFFFFFFF0;
    // rom_array[35918] = 32'hFFFFFFF0;
    // rom_array[35919] = 32'hFFFFFFF0;
    // rom_array[35920] = 32'hFFFFFFF0;
    // rom_array[35921] = 32'hFFFFFFF1;
    // rom_array[35922] = 32'hFFFFFFF1;
    // rom_array[35923] = 32'hFFFFFFF1;
    // rom_array[35924] = 32'hFFFFFFF1;
    // rom_array[35925] = 32'hFFFFFFF0;
    // rom_array[35926] = 32'hFFFFFFF0;
    // rom_array[35927] = 32'hFFFFFFF0;
    // rom_array[35928] = 32'hFFFFFFF0;
    // rom_array[35929] = 32'hFFFFFFF1;
    // rom_array[35930] = 32'hFFFFFFF1;
    // rom_array[35931] = 32'hFFFFFFF1;
    // rom_array[35932] = 32'hFFFFFFF1;
    // rom_array[35933] = 32'hFFFFFFF1;
    // rom_array[35934] = 32'hFFFFFFF1;
    // rom_array[35935] = 32'hFFFFFFF1;
    // rom_array[35936] = 32'hFFFFFFF1;
    // rom_array[35937] = 32'hFFFFFFF1;
    // rom_array[35938] = 32'hFFFFFFF1;
    // rom_array[35939] = 32'hFFFFFFF1;
    // rom_array[35940] = 32'hFFFFFFF1;
    // rom_array[35941] = 32'hFFFFFFF1;
    // rom_array[35942] = 32'hFFFFFFF1;
    // rom_array[35943] = 32'hFFFFFFF1;
    // rom_array[35944] = 32'hFFFFFFF1;
    // rom_array[35945] = 32'hFFFFFFF1;
    // rom_array[35946] = 32'hFFFFFFF1;
    // rom_array[35947] = 32'hFFFFFFF1;
    // rom_array[35948] = 32'hFFFFFFF1;
    // rom_array[35949] = 32'hFFFFFFF0;
    // rom_array[35950] = 32'hFFFFFFF0;
    // rom_array[35951] = 32'hFFFFFFF0;
    // rom_array[35952] = 32'hFFFFFFF0;
    // rom_array[35953] = 32'hFFFFFFF1;
    // rom_array[35954] = 32'hFFFFFFF1;
    // rom_array[35955] = 32'hFFFFFFF1;
    // rom_array[35956] = 32'hFFFFFFF1;
    // rom_array[35957] = 32'hFFFFFFF0;
    // rom_array[35958] = 32'hFFFFFFF0;
    // rom_array[35959] = 32'hFFFFFFF0;
    // rom_array[35960] = 32'hFFFFFFF0;
    // rom_array[35961] = 32'hFFFFFFF1;
    // rom_array[35962] = 32'hFFFFFFF1;
    // rom_array[35963] = 32'hFFFFFFF1;
    // rom_array[35964] = 32'hFFFFFFF1;
    // rom_array[35965] = 32'hFFFFFFF0;
    // rom_array[35966] = 32'hFFFFFFF0;
    // rom_array[35967] = 32'hFFFFFFF0;
    // rom_array[35968] = 32'hFFFFFFF0;
    // rom_array[35969] = 32'hFFFFFFF1;
    // rom_array[35970] = 32'hFFFFFFF1;
    // rom_array[35971] = 32'hFFFFFFF1;
    // rom_array[35972] = 32'hFFFFFFF1;
    // rom_array[35973] = 32'hFFFFFFF0;
    // rom_array[35974] = 32'hFFFFFFF0;
    // rom_array[35975] = 32'hFFFFFFF0;
    // rom_array[35976] = 32'hFFFFFFF0;
    // rom_array[35977] = 32'hFFFFFFF0;
    // rom_array[35978] = 32'hFFFFFFF0;
    // rom_array[35979] = 32'hFFFFFFF0;
    // rom_array[35980] = 32'hFFFFFFF0;
    // rom_array[35981] = 32'hFFFFFFF0;
    // rom_array[35982] = 32'hFFFFFFF0;
    // rom_array[35983] = 32'hFFFFFFF1;
    // rom_array[35984] = 32'hFFFFFFF1;
    // rom_array[35985] = 32'hFFFFFFF0;
    // rom_array[35986] = 32'hFFFFFFF0;
    // rom_array[35987] = 32'hFFFFFFF0;
    // rom_array[35988] = 32'hFFFFFFF0;
    // rom_array[35989] = 32'hFFFFFFF0;
    // rom_array[35990] = 32'hFFFFFFF0;
    // rom_array[35991] = 32'hFFFFFFF1;
    // rom_array[35992] = 32'hFFFFFFF1;
    // rom_array[35993] = 32'hFFFFFFF0;
    // rom_array[35994] = 32'hFFFFFFF0;
    // rom_array[35995] = 32'hFFFFFFF0;
    // rom_array[35996] = 32'hFFFFFFF0;
    // rom_array[35997] = 32'hFFFFFFF1;
    // rom_array[35998] = 32'hFFFFFFF1;
    // rom_array[35999] = 32'hFFFFFFF1;
    // rom_array[36000] = 32'hFFFFFFF1;
    // rom_array[36001] = 32'hFFFFFFF0;
    // rom_array[36002] = 32'hFFFFFFF0;
    // rom_array[36003] = 32'hFFFFFFF0;
    // rom_array[36004] = 32'hFFFFFFF0;
    // rom_array[36005] = 32'hFFFFFFF1;
    // rom_array[36006] = 32'hFFFFFFF1;
    // rom_array[36007] = 32'hFFFFFFF1;
    // rom_array[36008] = 32'hFFFFFFF1;
    // rom_array[36009] = 32'hFFFFFFF0;
    // rom_array[36010] = 32'hFFFFFFF0;
    // rom_array[36011] = 32'hFFFFFFF0;
    // rom_array[36012] = 32'hFFFFFFF0;
    // rom_array[36013] = 32'hFFFFFFF1;
    // rom_array[36014] = 32'hFFFFFFF1;
    // rom_array[36015] = 32'hFFFFFFF1;
    // rom_array[36016] = 32'hFFFFFFF1;
    // rom_array[36017] = 32'hFFFFFFF0;
    // rom_array[36018] = 32'hFFFFFFF0;
    // rom_array[36019] = 32'hFFFFFFF0;
    // rom_array[36020] = 32'hFFFFFFF0;
    // rom_array[36021] = 32'hFFFFFFF1;
    // rom_array[36022] = 32'hFFFFFFF1;
    // rom_array[36023] = 32'hFFFFFFF1;
    // rom_array[36024] = 32'hFFFFFFF1;
    // rom_array[36025] = 32'hFFFFFFF0;
    // rom_array[36026] = 32'hFFFFFFF0;
    // rom_array[36027] = 32'hFFFFFFF0;
    // rom_array[36028] = 32'hFFFFFFF0;
    // rom_array[36029] = 32'hFFFFFFF1;
    // rom_array[36030] = 32'hFFFFFFF1;
    // rom_array[36031] = 32'hFFFFFFF1;
    // rom_array[36032] = 32'hFFFFFFF1;
    // rom_array[36033] = 32'hFFFFFFF0;
    // rom_array[36034] = 32'hFFFFFFF0;
    // rom_array[36035] = 32'hFFFFFFF0;
    // rom_array[36036] = 32'hFFFFFFF0;
    // rom_array[36037] = 32'hFFFFFFF1;
    // rom_array[36038] = 32'hFFFFFFF1;
    // rom_array[36039] = 32'hFFFFFFF1;
    // rom_array[36040] = 32'hFFFFFFF1;
    // rom_array[36041] = 32'hFFFFFFF0;
    // rom_array[36042] = 32'hFFFFFFF0;
    // rom_array[36043] = 32'hFFFFFFF1;
    // rom_array[36044] = 32'hFFFFFFF1;
    // rom_array[36045] = 32'hFFFFFFF0;
    // rom_array[36046] = 32'hFFFFFFF0;
    // rom_array[36047] = 32'hFFFFFFF1;
    // rom_array[36048] = 32'hFFFFFFF1;
    // rom_array[36049] = 32'hFFFFFFF0;
    // rom_array[36050] = 32'hFFFFFFF0;
    // rom_array[36051] = 32'hFFFFFFF1;
    // rom_array[36052] = 32'hFFFFFFF1;
    // rom_array[36053] = 32'hFFFFFFF0;
    // rom_array[36054] = 32'hFFFFFFF0;
    // rom_array[36055] = 32'hFFFFFFF1;
    // rom_array[36056] = 32'hFFFFFFF1;
    // rom_array[36057] = 32'hFFFFFFF0;
    // rom_array[36058] = 32'hFFFFFFF0;
    // rom_array[36059] = 32'hFFFFFFF1;
    // rom_array[36060] = 32'hFFFFFFF1;
    // rom_array[36061] = 32'hFFFFFFF0;
    // rom_array[36062] = 32'hFFFFFFF0;
    // rom_array[36063] = 32'hFFFFFFF1;
    // rom_array[36064] = 32'hFFFFFFF1;
    // rom_array[36065] = 32'hFFFFFFF0;
    // rom_array[36066] = 32'hFFFFFFF0;
    // rom_array[36067] = 32'hFFFFFFF1;
    // rom_array[36068] = 32'hFFFFFFF1;
    // rom_array[36069] = 32'hFFFFFFF0;
    // rom_array[36070] = 32'hFFFFFFF0;
    // rom_array[36071] = 32'hFFFFFFF1;
    // rom_array[36072] = 32'hFFFFFFF1;
    // rom_array[36073] = 32'hFFFFFFF0;
    // rom_array[36074] = 32'hFFFFFFF0;
    // rom_array[36075] = 32'hFFFFFFF1;
    // rom_array[36076] = 32'hFFFFFFF1;
    // rom_array[36077] = 32'hFFFFFFF0;
    // rom_array[36078] = 32'hFFFFFFF0;
    // rom_array[36079] = 32'hFFFFFFF1;
    // rom_array[36080] = 32'hFFFFFFF1;
    // rom_array[36081] = 32'hFFFFFFF0;
    // rom_array[36082] = 32'hFFFFFFF0;
    // rom_array[36083] = 32'hFFFFFFF1;
    // rom_array[36084] = 32'hFFFFFFF1;
    // rom_array[36085] = 32'hFFFFFFF0;
    // rom_array[36086] = 32'hFFFFFFF0;
    // rom_array[36087] = 32'hFFFFFFF1;
    // rom_array[36088] = 32'hFFFFFFF1;
    // rom_array[36089] = 32'hFFFFFFF0;
    // rom_array[36090] = 32'hFFFFFFF0;
    // rom_array[36091] = 32'hFFFFFFF1;
    // rom_array[36092] = 32'hFFFFFFF1;
    // rom_array[36093] = 32'hFFFFFFF0;
    // rom_array[36094] = 32'hFFFFFFF0;
    // rom_array[36095] = 32'hFFFFFFF1;
    // rom_array[36096] = 32'hFFFFFFF1;
    // rom_array[36097] = 32'hFFFFFFF0;
    // rom_array[36098] = 32'hFFFFFFF0;
    // rom_array[36099] = 32'hFFFFFFF1;
    // rom_array[36100] = 32'hFFFFFFF1;
    // rom_array[36101] = 32'hFFFFFFF0;
    // rom_array[36102] = 32'hFFFFFFF0;
    // rom_array[36103] = 32'hFFFFFFF1;
    // rom_array[36104] = 32'hFFFFFFF1;
    // rom_array[36105] = 32'hFFFFFFF0;
    // rom_array[36106] = 32'hFFFFFFF0;
    // rom_array[36107] = 32'hFFFFFFF1;
    // rom_array[36108] = 32'hFFFFFFF1;
    // rom_array[36109] = 32'hFFFFFFF0;
    // rom_array[36110] = 32'hFFFFFFF0;
    // rom_array[36111] = 32'hFFFFFFF1;
    // rom_array[36112] = 32'hFFFFFFF1;
    // rom_array[36113] = 32'hFFFFFFF0;
    // rom_array[36114] = 32'hFFFFFFF0;
    // rom_array[36115] = 32'hFFFFFFF1;
    // rom_array[36116] = 32'hFFFFFFF1;
    // rom_array[36117] = 32'hFFFFFFF0;
    // rom_array[36118] = 32'hFFFFFFF0;
    // rom_array[36119] = 32'hFFFFFFF1;
    // rom_array[36120] = 32'hFFFFFFF1;
    // rom_array[36121] = 32'hFFFFFFF0;
    // rom_array[36122] = 32'hFFFFFFF0;
    // rom_array[36123] = 32'hFFFFFFF1;
    // rom_array[36124] = 32'hFFFFFFF1;
    // rom_array[36125] = 32'hFFFFFFF0;
    // rom_array[36126] = 32'hFFFFFFF0;
    // rom_array[36127] = 32'hFFFFFFF1;
    // rom_array[36128] = 32'hFFFFFFF1;
    // rom_array[36129] = 32'hFFFFFFF0;
    // rom_array[36130] = 32'hFFFFFFF0;
    // rom_array[36131] = 32'hFFFFFFF1;
    // rom_array[36132] = 32'hFFFFFFF1;
    // rom_array[36133] = 32'hFFFFFFF0;
    // rom_array[36134] = 32'hFFFFFFF0;
    // rom_array[36135] = 32'hFFFFFFF1;
    // rom_array[36136] = 32'hFFFFFFF1;
    // rom_array[36137] = 32'hFFFFFFF0;
    // rom_array[36138] = 32'hFFFFFFF0;
    // rom_array[36139] = 32'hFFFFFFF0;
    // rom_array[36140] = 32'hFFFFFFF0;
    // rom_array[36141] = 32'hFFFFFFF1;
    // rom_array[36142] = 32'hFFFFFFF1;
    // rom_array[36143] = 32'hFFFFFFF1;
    // rom_array[36144] = 32'hFFFFFFF1;
    // rom_array[36145] = 32'hFFFFFFF0;
    // rom_array[36146] = 32'hFFFFFFF0;
    // rom_array[36147] = 32'hFFFFFFF0;
    // rom_array[36148] = 32'hFFFFFFF0;
    // rom_array[36149] = 32'hFFFFFFF1;
    // rom_array[36150] = 32'hFFFFFFF1;
    // rom_array[36151] = 32'hFFFFFFF1;
    // rom_array[36152] = 32'hFFFFFFF1;
    // rom_array[36153] = 32'hFFFFFFF1;
    // rom_array[36154] = 32'hFFFFFFF1;
    // rom_array[36155] = 32'hFFFFFFF1;
    // rom_array[36156] = 32'hFFFFFFF1;
    // rom_array[36157] = 32'hFFFFFFF1;
    // rom_array[36158] = 32'hFFFFFFF1;
    // rom_array[36159] = 32'hFFFFFFF1;
    // rom_array[36160] = 32'hFFFFFFF1;
    // rom_array[36161] = 32'hFFFFFFF1;
    // rom_array[36162] = 32'hFFFFFFF1;
    // rom_array[36163] = 32'hFFFFFFF1;
    // rom_array[36164] = 32'hFFFFFFF1;
    // rom_array[36165] = 32'hFFFFFFF1;
    // rom_array[36166] = 32'hFFFFFFF1;
    // rom_array[36167] = 32'hFFFFFFF1;
    // rom_array[36168] = 32'hFFFFFFF1;
    // rom_array[36169] = 32'hFFFFFFF1;
    // rom_array[36170] = 32'hFFFFFFF1;
    // rom_array[36171] = 32'hFFFFFFF1;
    // rom_array[36172] = 32'hFFFFFFF1;
    // rom_array[36173] = 32'hFFFFFFF1;
    // rom_array[36174] = 32'hFFFFFFF1;
    // rom_array[36175] = 32'hFFFFFFF1;
    // rom_array[36176] = 32'hFFFFFFF1;
    // rom_array[36177] = 32'hFFFFFFF1;
    // rom_array[36178] = 32'hFFFFFFF1;
    // rom_array[36179] = 32'hFFFFFFF1;
    // rom_array[36180] = 32'hFFFFFFF1;
    // rom_array[36181] = 32'hFFFFFFF1;
    // rom_array[36182] = 32'hFFFFFFF1;
    // rom_array[36183] = 32'hFFFFFFF1;
    // rom_array[36184] = 32'hFFFFFFF1;
    // rom_array[36185] = 32'hFFFFFFF1;
    // rom_array[36186] = 32'hFFFFFFF1;
    // rom_array[36187] = 32'hFFFFFFF1;
    // rom_array[36188] = 32'hFFFFFFF1;
    // rom_array[36189] = 32'hFFFFFFF1;
    // rom_array[36190] = 32'hFFFFFFF1;
    // rom_array[36191] = 32'hFFFFFFF1;
    // rom_array[36192] = 32'hFFFFFFF1;
    // rom_array[36193] = 32'hFFFFFFF1;
    // rom_array[36194] = 32'hFFFFFFF1;
    // rom_array[36195] = 32'hFFFFFFF1;
    // rom_array[36196] = 32'hFFFFFFF1;
    // rom_array[36197] = 32'hFFFFFFF1;
    // rom_array[36198] = 32'hFFFFFFF1;
    // rom_array[36199] = 32'hFFFFFFF1;
    // rom_array[36200] = 32'hFFFFFFF1;
    // rom_array[36201] = 32'hFFFFFFF1;
    // rom_array[36202] = 32'hFFFFFFF1;
    // rom_array[36203] = 32'hFFFFFFF1;
    // rom_array[36204] = 32'hFFFFFFF1;
    // rom_array[36205] = 32'hFFFFFFF1;
    // rom_array[36206] = 32'hFFFFFFF1;
    // rom_array[36207] = 32'hFFFFFFF1;
    // rom_array[36208] = 32'hFFFFFFF1;
    // rom_array[36209] = 32'hFFFFFFF1;
    // rom_array[36210] = 32'hFFFFFFF1;
    // rom_array[36211] = 32'hFFFFFFF1;
    // rom_array[36212] = 32'hFFFFFFF1;
    // rom_array[36213] = 32'hFFFFFFF1;
    // rom_array[36214] = 32'hFFFFFFF1;
    // rom_array[36215] = 32'hFFFFFFF1;
    // rom_array[36216] = 32'hFFFFFFF1;
    // rom_array[36217] = 32'hFFFFFFF1;
    // rom_array[36218] = 32'hFFFFFFF1;
    // rom_array[36219] = 32'hFFFFFFF1;
    // rom_array[36220] = 32'hFFFFFFF1;
    // rom_array[36221] = 32'hFFFFFFF1;
    // rom_array[36222] = 32'hFFFFFFF1;
    // rom_array[36223] = 32'hFFFFFFF1;
    // rom_array[36224] = 32'hFFFFFFF1;
    // rom_array[36225] = 32'hFFFFFFF1;
    // rom_array[36226] = 32'hFFFFFFF1;
    // rom_array[36227] = 32'hFFFFFFF1;
    // rom_array[36228] = 32'hFFFFFFF1;
    // rom_array[36229] = 32'hFFFFFFF1;
    // rom_array[36230] = 32'hFFFFFFF1;
    // rom_array[36231] = 32'hFFFFFFF1;
    // rom_array[36232] = 32'hFFFFFFF1;
    // rom_array[36233] = 32'hFFFFFFF0;
    // rom_array[36234] = 32'hFFFFFFF0;
    // rom_array[36235] = 32'hFFFFFFF0;
    // rom_array[36236] = 32'hFFFFFFF0;
    // rom_array[36237] = 32'hFFFFFFF1;
    // rom_array[36238] = 32'hFFFFFFF1;
    // rom_array[36239] = 32'hFFFFFFF1;
    // rom_array[36240] = 32'hFFFFFFF1;
    // rom_array[36241] = 32'hFFFFFFF0;
    // rom_array[36242] = 32'hFFFFFFF0;
    // rom_array[36243] = 32'hFFFFFFF0;
    // rom_array[36244] = 32'hFFFFFFF0;
    // rom_array[36245] = 32'hFFFFFFF1;
    // rom_array[36246] = 32'hFFFFFFF1;
    // rom_array[36247] = 32'hFFFFFFF1;
    // rom_array[36248] = 32'hFFFFFFF1;
    // rom_array[36249] = 32'hFFFFFFF1;
    // rom_array[36250] = 32'hFFFFFFF1;
    // rom_array[36251] = 32'hFFFFFFF1;
    // rom_array[36252] = 32'hFFFFFFF1;
    // rom_array[36253] = 32'hFFFFFFF1;
    // rom_array[36254] = 32'hFFFFFFF1;
    // rom_array[36255] = 32'hFFFFFFF1;
    // rom_array[36256] = 32'hFFFFFFF1;
    // rom_array[36257] = 32'hFFFFFFF1;
    // rom_array[36258] = 32'hFFFFFFF1;
    // rom_array[36259] = 32'hFFFFFFF1;
    // rom_array[36260] = 32'hFFFFFFF1;
    // rom_array[36261] = 32'hFFFFFFF1;
    // rom_array[36262] = 32'hFFFFFFF1;
    // rom_array[36263] = 32'hFFFFFFF1;
    // rom_array[36264] = 32'hFFFFFFF1;
    // rom_array[36265] = 32'hFFFFFFF0;
    // rom_array[36266] = 32'hFFFFFFF0;
    // rom_array[36267] = 32'hFFFFFFF0;
    // rom_array[36268] = 32'hFFFFFFF0;
    // rom_array[36269] = 32'hFFFFFFF1;
    // rom_array[36270] = 32'hFFFFFFF1;
    // rom_array[36271] = 32'hFFFFFFF1;
    // rom_array[36272] = 32'hFFFFFFF1;
    // rom_array[36273] = 32'hFFFFFFF0;
    // rom_array[36274] = 32'hFFFFFFF0;
    // rom_array[36275] = 32'hFFFFFFF0;
    // rom_array[36276] = 32'hFFFFFFF0;
    // rom_array[36277] = 32'hFFFFFFF1;
    // rom_array[36278] = 32'hFFFFFFF1;
    // rom_array[36279] = 32'hFFFFFFF1;
    // rom_array[36280] = 32'hFFFFFFF1;
    // rom_array[36281] = 32'hFFFFFFF0;
    // rom_array[36282] = 32'hFFFFFFF0;
    // rom_array[36283] = 32'hFFFFFFF0;
    // rom_array[36284] = 32'hFFFFFFF0;
    // rom_array[36285] = 32'hFFFFFFF1;
    // rom_array[36286] = 32'hFFFFFFF1;
    // rom_array[36287] = 32'hFFFFFFF1;
    // rom_array[36288] = 32'hFFFFFFF1;
    // rom_array[36289] = 32'hFFFFFFF0;
    // rom_array[36290] = 32'hFFFFFFF0;
    // rom_array[36291] = 32'hFFFFFFF0;
    // rom_array[36292] = 32'hFFFFFFF0;
    // rom_array[36293] = 32'hFFFFFFF1;
    // rom_array[36294] = 32'hFFFFFFF1;
    // rom_array[36295] = 32'hFFFFFFF1;
    // rom_array[36296] = 32'hFFFFFFF1;
    // rom_array[36297] = 32'hFFFFFFF0;
    // rom_array[36298] = 32'hFFFFFFF0;
    // rom_array[36299] = 32'hFFFFFFF0;
    // rom_array[36300] = 32'hFFFFFFF0;
    // rom_array[36301] = 32'hFFFFFFF1;
    // rom_array[36302] = 32'hFFFFFFF1;
    // rom_array[36303] = 32'hFFFFFFF1;
    // rom_array[36304] = 32'hFFFFFFF1;
    // rom_array[36305] = 32'hFFFFFFF0;
    // rom_array[36306] = 32'hFFFFFFF0;
    // rom_array[36307] = 32'hFFFFFFF0;
    // rom_array[36308] = 32'hFFFFFFF0;
    // rom_array[36309] = 32'hFFFFFFF1;
    // rom_array[36310] = 32'hFFFFFFF1;
    // rom_array[36311] = 32'hFFFFFFF1;
    // rom_array[36312] = 32'hFFFFFFF1;
    // rom_array[36313] = 32'hFFFFFFF0;
    // rom_array[36314] = 32'hFFFFFFF0;
    // rom_array[36315] = 32'hFFFFFFF0;
    // rom_array[36316] = 32'hFFFFFFF0;
    // rom_array[36317] = 32'hFFFFFFF1;
    // rom_array[36318] = 32'hFFFFFFF1;
    // rom_array[36319] = 32'hFFFFFFF1;
    // rom_array[36320] = 32'hFFFFFFF1;
    // rom_array[36321] = 32'hFFFFFFF0;
    // rom_array[36322] = 32'hFFFFFFF0;
    // rom_array[36323] = 32'hFFFFFFF0;
    // rom_array[36324] = 32'hFFFFFFF0;
    // rom_array[36325] = 32'hFFFFFFF1;
    // rom_array[36326] = 32'hFFFFFFF1;
    // rom_array[36327] = 32'hFFFFFFF1;
    // rom_array[36328] = 32'hFFFFFFF1;
    // rom_array[36329] = 32'hFFFFFFF0;
    // rom_array[36330] = 32'hFFFFFFF0;
    // rom_array[36331] = 32'hFFFFFFF0;
    // rom_array[36332] = 32'hFFFFFFF0;
    // rom_array[36333] = 32'hFFFFFFF1;
    // rom_array[36334] = 32'hFFFFFFF1;
    // rom_array[36335] = 32'hFFFFFFF1;
    // rom_array[36336] = 32'hFFFFFFF1;
    // rom_array[36337] = 32'hFFFFFFF0;
    // rom_array[36338] = 32'hFFFFFFF0;
    // rom_array[36339] = 32'hFFFFFFF0;
    // rom_array[36340] = 32'hFFFFFFF0;
    // rom_array[36341] = 32'hFFFFFFF1;
    // rom_array[36342] = 32'hFFFFFFF1;
    // rom_array[36343] = 32'hFFFFFFF1;
    // rom_array[36344] = 32'hFFFFFFF1;
    // rom_array[36345] = 32'hFFFFFFF0;
    // rom_array[36346] = 32'hFFFFFFF0;
    // rom_array[36347] = 32'hFFFFFFF0;
    // rom_array[36348] = 32'hFFFFFFF0;
    // rom_array[36349] = 32'hFFFFFFF1;
    // rom_array[36350] = 32'hFFFFFFF1;
    // rom_array[36351] = 32'hFFFFFFF1;
    // rom_array[36352] = 32'hFFFFFFF1;
    // rom_array[36353] = 32'hFFFFFFF0;
    // rom_array[36354] = 32'hFFFFFFF0;
    // rom_array[36355] = 32'hFFFFFFF0;
    // rom_array[36356] = 32'hFFFFFFF0;
    // rom_array[36357] = 32'hFFFFFFF1;
    // rom_array[36358] = 32'hFFFFFFF1;
    // rom_array[36359] = 32'hFFFFFFF1;
    // rom_array[36360] = 32'hFFFFFFF1;
    // rom_array[36361] = 32'hFFFFFFF0;
    // rom_array[36362] = 32'hFFFFFFF0;
    // rom_array[36363] = 32'hFFFFFFF1;
    // rom_array[36364] = 32'hFFFFFFF1;
    // rom_array[36365] = 32'hFFFFFFF0;
    // rom_array[36366] = 32'hFFFFFFF0;
    // rom_array[36367] = 32'hFFFFFFF1;
    // rom_array[36368] = 32'hFFFFFFF1;
    // rom_array[36369] = 32'hFFFFFFF0;
    // rom_array[36370] = 32'hFFFFFFF0;
    // rom_array[36371] = 32'hFFFFFFF1;
    // rom_array[36372] = 32'hFFFFFFF1;
    // rom_array[36373] = 32'hFFFFFFF0;
    // rom_array[36374] = 32'hFFFFFFF0;
    // rom_array[36375] = 32'hFFFFFFF1;
    // rom_array[36376] = 32'hFFFFFFF1;
    // rom_array[36377] = 32'hFFFFFFF0;
    // rom_array[36378] = 32'hFFFFFFF0;
    // rom_array[36379] = 32'hFFFFFFF1;
    // rom_array[36380] = 32'hFFFFFFF1;
    // rom_array[36381] = 32'hFFFFFFF0;
    // rom_array[36382] = 32'hFFFFFFF0;
    // rom_array[36383] = 32'hFFFFFFF1;
    // rom_array[36384] = 32'hFFFFFFF1;
    // rom_array[36385] = 32'hFFFFFFF0;
    // rom_array[36386] = 32'hFFFFFFF0;
    // rom_array[36387] = 32'hFFFFFFF1;
    // rom_array[36388] = 32'hFFFFFFF1;
    // rom_array[36389] = 32'hFFFFFFF0;
    // rom_array[36390] = 32'hFFFFFFF0;
    // rom_array[36391] = 32'hFFFFFFF1;
    // rom_array[36392] = 32'hFFFFFFF1;
    // rom_array[36393] = 32'hFFFFFFF0;
    // rom_array[36394] = 32'hFFFFFFF0;
    // rom_array[36395] = 32'hFFFFFFF1;
    // rom_array[36396] = 32'hFFFFFFF1;
    // rom_array[36397] = 32'hFFFFFFF0;
    // rom_array[36398] = 32'hFFFFFFF0;
    // rom_array[36399] = 32'hFFFFFFF1;
    // rom_array[36400] = 32'hFFFFFFF1;
    // rom_array[36401] = 32'hFFFFFFF0;
    // rom_array[36402] = 32'hFFFFFFF0;
    // rom_array[36403] = 32'hFFFFFFF1;
    // rom_array[36404] = 32'hFFFFFFF1;
    // rom_array[36405] = 32'hFFFFFFF0;
    // rom_array[36406] = 32'hFFFFFFF0;
    // rom_array[36407] = 32'hFFFFFFF1;
    // rom_array[36408] = 32'hFFFFFFF1;
    // rom_array[36409] = 32'hFFFFFFF0;
    // rom_array[36410] = 32'hFFFFFFF0;
    // rom_array[36411] = 32'hFFFFFFF1;
    // rom_array[36412] = 32'hFFFFFFF1;
    // rom_array[36413] = 32'hFFFFFFF0;
    // rom_array[36414] = 32'hFFFFFFF0;
    // rom_array[36415] = 32'hFFFFFFF1;
    // rom_array[36416] = 32'hFFFFFFF1;
    // rom_array[36417] = 32'hFFFFFFF0;
    // rom_array[36418] = 32'hFFFFFFF0;
    // rom_array[36419] = 32'hFFFFFFF1;
    // rom_array[36420] = 32'hFFFFFFF1;
    // rom_array[36421] = 32'hFFFFFFF0;
    // rom_array[36422] = 32'hFFFFFFF0;
    // rom_array[36423] = 32'hFFFFFFF1;
    // rom_array[36424] = 32'hFFFFFFF1;
    // rom_array[36425] = 32'hFFFFFFF0;
    // rom_array[36426] = 32'hFFFFFFF0;
    // rom_array[36427] = 32'hFFFFFFF1;
    // rom_array[36428] = 32'hFFFFFFF1;
    // rom_array[36429] = 32'hFFFFFFF0;
    // rom_array[36430] = 32'hFFFFFFF0;
    // rom_array[36431] = 32'hFFFFFFF1;
    // rom_array[36432] = 32'hFFFFFFF1;
    // rom_array[36433] = 32'hFFFFFFF0;
    // rom_array[36434] = 32'hFFFFFFF0;
    // rom_array[36435] = 32'hFFFFFFF1;
    // rom_array[36436] = 32'hFFFFFFF1;
    // rom_array[36437] = 32'hFFFFFFF0;
    // rom_array[36438] = 32'hFFFFFFF0;
    // rom_array[36439] = 32'hFFFFFFF1;
    // rom_array[36440] = 32'hFFFFFFF1;
    // rom_array[36441] = 32'hFFFFFFF0;
    // rom_array[36442] = 32'hFFFFFFF0;
    // rom_array[36443] = 32'hFFFFFFF1;
    // rom_array[36444] = 32'hFFFFFFF1;
    // rom_array[36445] = 32'hFFFFFFF0;
    // rom_array[36446] = 32'hFFFFFFF0;
    // rom_array[36447] = 32'hFFFFFFF1;
    // rom_array[36448] = 32'hFFFFFFF1;
    // rom_array[36449] = 32'hFFFFFFF0;
    // rom_array[36450] = 32'hFFFFFFF0;
    // rom_array[36451] = 32'hFFFFFFF1;
    // rom_array[36452] = 32'hFFFFFFF1;
    // rom_array[36453] = 32'hFFFFFFF0;
    // rom_array[36454] = 32'hFFFFFFF0;
    // rom_array[36455] = 32'hFFFFFFF1;
    // rom_array[36456] = 32'hFFFFFFF1;
    // rom_array[36457] = 32'hFFFFFFF0;
    // rom_array[36458] = 32'hFFFFFFF0;
    // rom_array[36459] = 32'hFFFFFFF1;
    // rom_array[36460] = 32'hFFFFFFF1;
    // rom_array[36461] = 32'hFFFFFFF0;
    // rom_array[36462] = 32'hFFFFFFF0;
    // rom_array[36463] = 32'hFFFFFFF1;
    // rom_array[36464] = 32'hFFFFFFF1;
    // rom_array[36465] = 32'hFFFFFFF0;
    // rom_array[36466] = 32'hFFFFFFF0;
    // rom_array[36467] = 32'hFFFFFFF1;
    // rom_array[36468] = 32'hFFFFFFF1;
    // rom_array[36469] = 32'hFFFFFFF0;
    // rom_array[36470] = 32'hFFFFFFF0;
    // rom_array[36471] = 32'hFFFFFFF1;
    // rom_array[36472] = 32'hFFFFFFF1;
    // rom_array[36473] = 32'hFFFFFFF0;
    // rom_array[36474] = 32'hFFFFFFF0;
    // rom_array[36475] = 32'hFFFFFFF1;
    // rom_array[36476] = 32'hFFFFFFF1;
    // rom_array[36477] = 32'hFFFFFFF0;
    // rom_array[36478] = 32'hFFFFFFF0;
    // rom_array[36479] = 32'hFFFFFFF0;
    // rom_array[36480] = 32'hFFFFFFF0;
    // rom_array[36481] = 32'hFFFFFFF0;
    // rom_array[36482] = 32'hFFFFFFF0;
    // rom_array[36483] = 32'hFFFFFFF1;
    // rom_array[36484] = 32'hFFFFFFF1;
    // rom_array[36485] = 32'hFFFFFFF0;
    // rom_array[36486] = 32'hFFFFFFF0;
    // rom_array[36487] = 32'hFFFFFFF0;
    // rom_array[36488] = 32'hFFFFFFF0;
    // rom_array[36489] = 32'hFFFFFFF1;
    // rom_array[36490] = 32'hFFFFFFF1;
    // rom_array[36491] = 32'hFFFFFFF1;
    // rom_array[36492] = 32'hFFFFFFF1;
    // rom_array[36493] = 32'hFFFFFFF0;
    // rom_array[36494] = 32'hFFFFFFF0;
    // rom_array[36495] = 32'hFFFFFFF0;
    // rom_array[36496] = 32'hFFFFFFF0;
    // rom_array[36497] = 32'hFFFFFFF1;
    // rom_array[36498] = 32'hFFFFFFF1;
    // rom_array[36499] = 32'hFFFFFFF1;
    // rom_array[36500] = 32'hFFFFFFF1;
    // rom_array[36501] = 32'hFFFFFFF0;
    // rom_array[36502] = 32'hFFFFFFF0;
    // rom_array[36503] = 32'hFFFFFFF0;
    // rom_array[36504] = 32'hFFFFFFF0;
    // rom_array[36505] = 32'hFFFFFFF1;
    // rom_array[36506] = 32'hFFFFFFF1;
    // rom_array[36507] = 32'hFFFFFFF1;
    // rom_array[36508] = 32'hFFFFFFF1;
    // rom_array[36509] = 32'hFFFFFFF0;
    // rom_array[36510] = 32'hFFFFFFF0;
    // rom_array[36511] = 32'hFFFFFFF0;
    // rom_array[36512] = 32'hFFFFFFF0;
    // rom_array[36513] = 32'hFFFFFFF1;
    // rom_array[36514] = 32'hFFFFFFF1;
    // rom_array[36515] = 32'hFFFFFFF1;
    // rom_array[36516] = 32'hFFFFFFF1;
    // rom_array[36517] = 32'hFFFFFFF0;
    // rom_array[36518] = 32'hFFFFFFF0;
    // rom_array[36519] = 32'hFFFFFFF0;
    // rom_array[36520] = 32'hFFFFFFF0;
    // rom_array[36521] = 32'hFFFFFFF1;
    // rom_array[36522] = 32'hFFFFFFF1;
    // rom_array[36523] = 32'hFFFFFFF1;
    // rom_array[36524] = 32'hFFFFFFF1;
    // rom_array[36525] = 32'hFFFFFFF0;
    // rom_array[36526] = 32'hFFFFFFF0;
    // rom_array[36527] = 32'hFFFFFFF0;
    // rom_array[36528] = 32'hFFFFFFF0;
    // rom_array[36529] = 32'hFFFFFFF1;
    // rom_array[36530] = 32'hFFFFFFF1;
    // rom_array[36531] = 32'hFFFFFFF1;
    // rom_array[36532] = 32'hFFFFFFF1;
    // rom_array[36533] = 32'hFFFFFFF0;
    // rom_array[36534] = 32'hFFFFFFF0;
    // rom_array[36535] = 32'hFFFFFFF0;
    // rom_array[36536] = 32'hFFFFFFF0;
    // rom_array[36537] = 32'hFFFFFFF1;
    // rom_array[36538] = 32'hFFFFFFF1;
    // rom_array[36539] = 32'hFFFFFFF1;
    // rom_array[36540] = 32'hFFFFFFF1;
    // rom_array[36541] = 32'hFFFFFFF1;
    // rom_array[36542] = 32'hFFFFFFF1;
    // rom_array[36543] = 32'hFFFFFFF1;
    // rom_array[36544] = 32'hFFFFFFF1;
    // rom_array[36545] = 32'hFFFFFFF1;
    // rom_array[36546] = 32'hFFFFFFF1;
    // rom_array[36547] = 32'hFFFFFFF1;
    // rom_array[36548] = 32'hFFFFFFF1;
    // rom_array[36549] = 32'hFFFFFFF1;
    // rom_array[36550] = 32'hFFFFFFF1;
    // rom_array[36551] = 32'hFFFFFFF1;
    // rom_array[36552] = 32'hFFFFFFF1;
    // rom_array[36553] = 32'hFFFFFFF1;
    // rom_array[36554] = 32'hFFFFFFF1;
    // rom_array[36555] = 32'hFFFFFFF1;
    // rom_array[36556] = 32'hFFFFFFF1;
    // rom_array[36557] = 32'hFFFFFFF1;
    // rom_array[36558] = 32'hFFFFFFF1;
    // rom_array[36559] = 32'hFFFFFFF1;
    // rom_array[36560] = 32'hFFFFFFF1;
    // rom_array[36561] = 32'hFFFFFFF1;
    // rom_array[36562] = 32'hFFFFFFF1;
    // rom_array[36563] = 32'hFFFFFFF1;
    // rom_array[36564] = 32'hFFFFFFF1;
    // rom_array[36565] = 32'hFFFFFFF1;
    // rom_array[36566] = 32'hFFFFFFF1;
    // rom_array[36567] = 32'hFFFFFFF1;
    // rom_array[36568] = 32'hFFFFFFF1;
    // rom_array[36569] = 32'hFFFFFFF1;
    // rom_array[36570] = 32'hFFFFFFF1;
    // rom_array[36571] = 32'hFFFFFFF1;
    // rom_array[36572] = 32'hFFFFFFF1;
    // rom_array[36573] = 32'hFFFFFFF1;
    // rom_array[36574] = 32'hFFFFFFF1;
    // rom_array[36575] = 32'hFFFFFFF1;
    // rom_array[36576] = 32'hFFFFFFF1;
    // rom_array[36577] = 32'hFFFFFFF1;
    // rom_array[36578] = 32'hFFFFFFF1;
    // rom_array[36579] = 32'hFFFFFFF1;
    // rom_array[36580] = 32'hFFFFFFF1;
    // rom_array[36581] = 32'hFFFFFFF1;
    // rom_array[36582] = 32'hFFFFFFF1;
    // rom_array[36583] = 32'hFFFFFFF1;
    // rom_array[36584] = 32'hFFFFFFF1;
    // rom_array[36585] = 32'hFFFFFFF1;
    // rom_array[36586] = 32'hFFFFFFF1;
    // rom_array[36587] = 32'hFFFFFFF1;
    // rom_array[36588] = 32'hFFFFFFF1;
    // rom_array[36589] = 32'hFFFFFFF0;
    // rom_array[36590] = 32'hFFFFFFF0;
    // rom_array[36591] = 32'hFFFFFFF0;
    // rom_array[36592] = 32'hFFFFFFF0;
    // rom_array[36593] = 32'hFFFFFFF1;
    // rom_array[36594] = 32'hFFFFFFF1;
    // rom_array[36595] = 32'hFFFFFFF1;
    // rom_array[36596] = 32'hFFFFFFF1;
    // rom_array[36597] = 32'hFFFFFFF0;
    // rom_array[36598] = 32'hFFFFFFF0;
    // rom_array[36599] = 32'hFFFFFFF0;
    // rom_array[36600] = 32'hFFFFFFF0;
    // rom_array[36601] = 32'hFFFFFFF1;
    // rom_array[36602] = 32'hFFFFFFF1;
    // rom_array[36603] = 32'hFFFFFFF1;
    // rom_array[36604] = 32'hFFFFFFF1;
    // rom_array[36605] = 32'hFFFFFFF1;
    // rom_array[36606] = 32'hFFFFFFF1;
    // rom_array[36607] = 32'hFFFFFFF1;
    // rom_array[36608] = 32'hFFFFFFF1;
    // rom_array[36609] = 32'hFFFFFFF1;
    // rom_array[36610] = 32'hFFFFFFF1;
    // rom_array[36611] = 32'hFFFFFFF1;
    // rom_array[36612] = 32'hFFFFFFF1;
    // rom_array[36613] = 32'hFFFFFFF1;
    // rom_array[36614] = 32'hFFFFFFF1;
    // rom_array[36615] = 32'hFFFFFFF1;
    // rom_array[36616] = 32'hFFFFFFF1;
    // rom_array[36617] = 32'hFFFFFFF1;
    // rom_array[36618] = 32'hFFFFFFF1;
    // rom_array[36619] = 32'hFFFFFFF1;
    // rom_array[36620] = 32'hFFFFFFF1;
    // rom_array[36621] = 32'hFFFFFFF0;
    // rom_array[36622] = 32'hFFFFFFF0;
    // rom_array[36623] = 32'hFFFFFFF0;
    // rom_array[36624] = 32'hFFFFFFF0;
    // rom_array[36625] = 32'hFFFFFFF1;
    // rom_array[36626] = 32'hFFFFFFF1;
    // rom_array[36627] = 32'hFFFFFFF1;
    // rom_array[36628] = 32'hFFFFFFF1;
    // rom_array[36629] = 32'hFFFFFFF0;
    // rom_array[36630] = 32'hFFFFFFF0;
    // rom_array[36631] = 32'hFFFFFFF0;
    // rom_array[36632] = 32'hFFFFFFF0;
    // rom_array[36633] = 32'hFFFFFFF1;
    // rom_array[36634] = 32'hFFFFFFF1;
    // rom_array[36635] = 32'hFFFFFFF1;
    // rom_array[36636] = 32'hFFFFFFF1;
    // rom_array[36637] = 32'hFFFFFFF0;
    // rom_array[36638] = 32'hFFFFFFF0;
    // rom_array[36639] = 32'hFFFFFFF0;
    // rom_array[36640] = 32'hFFFFFFF0;
    // rom_array[36641] = 32'hFFFFFFF1;
    // rom_array[36642] = 32'hFFFFFFF1;
    // rom_array[36643] = 32'hFFFFFFF1;
    // rom_array[36644] = 32'hFFFFFFF1;
    // rom_array[36645] = 32'hFFFFFFF0;
    // rom_array[36646] = 32'hFFFFFFF0;
    // rom_array[36647] = 32'hFFFFFFF0;
    // rom_array[36648] = 32'hFFFFFFF0;
    // rom_array[36649] = 32'hFFFFFFF1;
    // rom_array[36650] = 32'hFFFFFFF1;
    // rom_array[36651] = 32'hFFFFFFF1;
    // rom_array[36652] = 32'hFFFFFFF1;
    // rom_array[36653] = 32'hFFFFFFF0;
    // rom_array[36654] = 32'hFFFFFFF0;
    // rom_array[36655] = 32'hFFFFFFF0;
    // rom_array[36656] = 32'hFFFFFFF0;
    // rom_array[36657] = 32'hFFFFFFF1;
    // rom_array[36658] = 32'hFFFFFFF1;
    // rom_array[36659] = 32'hFFFFFFF1;
    // rom_array[36660] = 32'hFFFFFFF1;
    // rom_array[36661] = 32'hFFFFFFF0;
    // rom_array[36662] = 32'hFFFFFFF0;
    // rom_array[36663] = 32'hFFFFFFF0;
    // rom_array[36664] = 32'hFFFFFFF0;
    // rom_array[36665] = 32'hFFFFFFF1;
    // rom_array[36666] = 32'hFFFFFFF1;
    // rom_array[36667] = 32'hFFFFFFF1;
    // rom_array[36668] = 32'hFFFFFFF1;
    // rom_array[36669] = 32'hFFFFFFF0;
    // rom_array[36670] = 32'hFFFFFFF0;
    // rom_array[36671] = 32'hFFFFFFF0;
    // rom_array[36672] = 32'hFFFFFFF0;
    // rom_array[36673] = 32'hFFFFFFF1;
    // rom_array[36674] = 32'hFFFFFFF1;
    // rom_array[36675] = 32'hFFFFFFF1;
    // rom_array[36676] = 32'hFFFFFFF1;
    // rom_array[36677] = 32'hFFFFFFF0;
    // rom_array[36678] = 32'hFFFFFFF0;
    // rom_array[36679] = 32'hFFFFFFF0;
    // rom_array[36680] = 32'hFFFFFFF0;
    // rom_array[36681] = 32'hFFFFFFF1;
    // rom_array[36682] = 32'hFFFFFFF1;
    // rom_array[36683] = 32'hFFFFFFF1;
    // rom_array[36684] = 32'hFFFFFFF1;
    // rom_array[36685] = 32'hFFFFFFF0;
    // rom_array[36686] = 32'hFFFFFFF0;
    // rom_array[36687] = 32'hFFFFFFF0;
    // rom_array[36688] = 32'hFFFFFFF0;
    // rom_array[36689] = 32'hFFFFFFF1;
    // rom_array[36690] = 32'hFFFFFFF1;
    // rom_array[36691] = 32'hFFFFFFF1;
    // rom_array[36692] = 32'hFFFFFFF1;
    // rom_array[36693] = 32'hFFFFFFF0;
    // rom_array[36694] = 32'hFFFFFFF0;
    // rom_array[36695] = 32'hFFFFFFF0;
    // rom_array[36696] = 32'hFFFFFFF0;
    // rom_array[36697] = 32'hFFFFFFF1;
    // rom_array[36698] = 32'hFFFFFFF1;
    // rom_array[36699] = 32'hFFFFFFF1;
    // rom_array[36700] = 32'hFFFFFFF1;
    // rom_array[36701] = 32'hFFFFFFF0;
    // rom_array[36702] = 32'hFFFFFFF0;
    // rom_array[36703] = 32'hFFFFFFF0;
    // rom_array[36704] = 32'hFFFFFFF0;
    // rom_array[36705] = 32'hFFFFFFF1;
    // rom_array[36706] = 32'hFFFFFFF1;
    // rom_array[36707] = 32'hFFFFFFF1;
    // rom_array[36708] = 32'hFFFFFFF1;
    // rom_array[36709] = 32'hFFFFFFF0;
    // rom_array[36710] = 32'hFFFFFFF0;
    // rom_array[36711] = 32'hFFFFFFF0;
    // rom_array[36712] = 32'hFFFFFFF0;
    // rom_array[36713] = 32'hFFFFFFF1;
    // rom_array[36714] = 32'hFFFFFFF1;
    // rom_array[36715] = 32'hFFFFFFF1;
    // rom_array[36716] = 32'hFFFFFFF1;
    // rom_array[36717] = 32'hFFFFFFF1;
    // rom_array[36718] = 32'hFFFFFFF1;
    // rom_array[36719] = 32'hFFFFFFF1;
    // rom_array[36720] = 32'hFFFFFFF1;
    // rom_array[36721] = 32'hFFFFFFF1;
    // rom_array[36722] = 32'hFFFFFFF1;
    // rom_array[36723] = 32'hFFFFFFF1;
    // rom_array[36724] = 32'hFFFFFFF1;
    // rom_array[36725] = 32'hFFFFFFF1;
    // rom_array[36726] = 32'hFFFFFFF1;
    // rom_array[36727] = 32'hFFFFFFF1;
    // rom_array[36728] = 32'hFFFFFFF1;
    // rom_array[36729] = 32'hFFFFFFF1;
    // rom_array[36730] = 32'hFFFFFFF1;
    // rom_array[36731] = 32'hFFFFFFF1;
    // rom_array[36732] = 32'hFFFFFFF1;
    // rom_array[36733] = 32'hFFFFFFF1;
    // rom_array[36734] = 32'hFFFFFFF1;
    // rom_array[36735] = 32'hFFFFFFF1;
    // rom_array[36736] = 32'hFFFFFFF1;
    // rom_array[36737] = 32'hFFFFFFF1;
    // rom_array[36738] = 32'hFFFFFFF1;
    // rom_array[36739] = 32'hFFFFFFF1;
    // rom_array[36740] = 32'hFFFFFFF1;
    // rom_array[36741] = 32'hFFFFFFF1;
    // rom_array[36742] = 32'hFFFFFFF1;
    // rom_array[36743] = 32'hFFFFFFF1;
    // rom_array[36744] = 32'hFFFFFFF1;
    // rom_array[36745] = 32'hFFFFFFF1;
    // rom_array[36746] = 32'hFFFFFFF1;
    // rom_array[36747] = 32'hFFFFFFF1;
    // rom_array[36748] = 32'hFFFFFFF1;
    // rom_array[36749] = 32'hFFFFFFF1;
    // rom_array[36750] = 32'hFFFFFFF1;
    // rom_array[36751] = 32'hFFFFFFF1;
    // rom_array[36752] = 32'hFFFFFFF1;
    // rom_array[36753] = 32'hFFFFFFF1;
    // rom_array[36754] = 32'hFFFFFFF1;
    // rom_array[36755] = 32'hFFFFFFF1;
    // rom_array[36756] = 32'hFFFFFFF1;
    // rom_array[36757] = 32'hFFFFFFF1;
    // rom_array[36758] = 32'hFFFFFFF1;
    // rom_array[36759] = 32'hFFFFFFF1;
    // rom_array[36760] = 32'hFFFFFFF1;
    // rom_array[36761] = 32'hFFFFFFF1;
    // rom_array[36762] = 32'hFFFFFFF1;
    // rom_array[36763] = 32'hFFFFFFF1;
    // rom_array[36764] = 32'hFFFFFFF1;
    // rom_array[36765] = 32'hFFFFFFF0;
    // rom_array[36766] = 32'hFFFFFFF0;
    // rom_array[36767] = 32'hFFFFFFF0;
    // rom_array[36768] = 32'hFFFFFFF0;
    // rom_array[36769] = 32'hFFFFFFF1;
    // rom_array[36770] = 32'hFFFFFFF1;
    // rom_array[36771] = 32'hFFFFFFF1;
    // rom_array[36772] = 32'hFFFFFFF1;
    // rom_array[36773] = 32'hFFFFFFF0;
    // rom_array[36774] = 32'hFFFFFFF0;
    // rom_array[36775] = 32'hFFFFFFF0;
    // rom_array[36776] = 32'hFFFFFFF0;
    // rom_array[36777] = 32'hFFFFFFF0;
    // rom_array[36778] = 32'hFFFFFFF0;
    // rom_array[36779] = 32'hFFFFFFF0;
    // rom_array[36780] = 32'hFFFFFFF0;
    // rom_array[36781] = 32'hFFFFFFF0;
    // rom_array[36782] = 32'hFFFFFFF0;
    // rom_array[36783] = 32'hFFFFFFF1;
    // rom_array[36784] = 32'hFFFFFFF1;
    // rom_array[36785] = 32'hFFFFFFF0;
    // rom_array[36786] = 32'hFFFFFFF0;
    // rom_array[36787] = 32'hFFFFFFF0;
    // rom_array[36788] = 32'hFFFFFFF0;
    // rom_array[36789] = 32'hFFFFFFF0;
    // rom_array[36790] = 32'hFFFFFFF0;
    // rom_array[36791] = 32'hFFFFFFF1;
    // rom_array[36792] = 32'hFFFFFFF1;
    // rom_array[36793] = 32'hFFFFFFF0;
    // rom_array[36794] = 32'hFFFFFFF0;
    // rom_array[36795] = 32'hFFFFFFF0;
    // rom_array[36796] = 32'hFFFFFFF0;
    // rom_array[36797] = 32'hFFFFFFF1;
    // rom_array[36798] = 32'hFFFFFFF1;
    // rom_array[36799] = 32'hFFFFFFF1;
    // rom_array[36800] = 32'hFFFFFFF1;
    // rom_array[36801] = 32'hFFFFFFF0;
    // rom_array[36802] = 32'hFFFFFFF0;
    // rom_array[36803] = 32'hFFFFFFF0;
    // rom_array[36804] = 32'hFFFFFFF0;
    // rom_array[36805] = 32'hFFFFFFF1;
    // rom_array[36806] = 32'hFFFFFFF1;
    // rom_array[36807] = 32'hFFFFFFF1;
    // rom_array[36808] = 32'hFFFFFFF1;
    // rom_array[36809] = 32'hFFFFFFF0;
    // rom_array[36810] = 32'hFFFFFFF0;
    // rom_array[36811] = 32'hFFFFFFF1;
    // rom_array[36812] = 32'hFFFFFFF1;
    // rom_array[36813] = 32'hFFFFFFF0;
    // rom_array[36814] = 32'hFFFFFFF0;
    // rom_array[36815] = 32'hFFFFFFF1;
    // rom_array[36816] = 32'hFFFFFFF1;
    // rom_array[36817] = 32'hFFFFFFF0;
    // rom_array[36818] = 32'hFFFFFFF0;
    // rom_array[36819] = 32'hFFFFFFF1;
    // rom_array[36820] = 32'hFFFFFFF1;
    // rom_array[36821] = 32'hFFFFFFF0;
    // rom_array[36822] = 32'hFFFFFFF0;
    // rom_array[36823] = 32'hFFFFFFF1;
    // rom_array[36824] = 32'hFFFFFFF1;
    // rom_array[36825] = 32'hFFFFFFF0;
    // rom_array[36826] = 32'hFFFFFFF0;
    // rom_array[36827] = 32'hFFFFFFF0;
    // rom_array[36828] = 32'hFFFFFFF0;
    // rom_array[36829] = 32'hFFFFFFF1;
    // rom_array[36830] = 32'hFFFFFFF1;
    // rom_array[36831] = 32'hFFFFFFF1;
    // rom_array[36832] = 32'hFFFFFFF1;
    // rom_array[36833] = 32'hFFFFFFF0;
    // rom_array[36834] = 32'hFFFFFFF0;
    // rom_array[36835] = 32'hFFFFFFF0;
    // rom_array[36836] = 32'hFFFFFFF0;
    // rom_array[36837] = 32'hFFFFFFF1;
    // rom_array[36838] = 32'hFFFFFFF1;
    // rom_array[36839] = 32'hFFFFFFF1;
    // rom_array[36840] = 32'hFFFFFFF1;
    // rom_array[36841] = 32'hFFFFFFF0;
    // rom_array[36842] = 32'hFFFFFFF0;
    // rom_array[36843] = 32'hFFFFFFF0;
    // rom_array[36844] = 32'hFFFFFFF0;
    // rom_array[36845] = 32'hFFFFFFF1;
    // rom_array[36846] = 32'hFFFFFFF1;
    // rom_array[36847] = 32'hFFFFFFF1;
    // rom_array[36848] = 32'hFFFFFFF1;
    // rom_array[36849] = 32'hFFFFFFF0;
    // rom_array[36850] = 32'hFFFFFFF0;
    // rom_array[36851] = 32'hFFFFFFF0;
    // rom_array[36852] = 32'hFFFFFFF0;
    // rom_array[36853] = 32'hFFFFFFF1;
    // rom_array[36854] = 32'hFFFFFFF1;
    // rom_array[36855] = 32'hFFFFFFF1;
    // rom_array[36856] = 32'hFFFFFFF1;
    // rom_array[36857] = 32'hFFFFFFF0;
    // rom_array[36858] = 32'hFFFFFFF0;
    // rom_array[36859] = 32'hFFFFFFF0;
    // rom_array[36860] = 32'hFFFFFFF0;
    // rom_array[36861] = 32'hFFFFFFF1;
    // rom_array[36862] = 32'hFFFFFFF1;
    // rom_array[36863] = 32'hFFFFFFF1;
    // rom_array[36864] = 32'hFFFFFFF1;
    // rom_array[36865] = 32'hFFFFFFF0;
    // rom_array[36866] = 32'hFFFFFFF0;
    // rom_array[36867] = 32'hFFFFFFF0;
    // rom_array[36868] = 32'hFFFFFFF0;
    // rom_array[36869] = 32'hFFFFFFF1;
    // rom_array[36870] = 32'hFFFFFFF1;
    // rom_array[36871] = 32'hFFFFFFF1;
    // rom_array[36872] = 32'hFFFFFFF1;
    // rom_array[36873] = 32'hFFFFFFF1;
    // rom_array[36874] = 32'hFFFFFFF1;
    // rom_array[36875] = 32'hFFFFFFF0;
    // rom_array[36876] = 32'hFFFFFFF0;
    // rom_array[36877] = 32'hFFFFFFF1;
    // rom_array[36878] = 32'hFFFFFFF1;
    // rom_array[36879] = 32'hFFFFFFF1;
    // rom_array[36880] = 32'hFFFFFFF1;
    // rom_array[36881] = 32'hFFFFFFF1;
    // rom_array[36882] = 32'hFFFFFFF1;
    // rom_array[36883] = 32'hFFFFFFF0;
    // rom_array[36884] = 32'hFFFFFFF0;
    // rom_array[36885] = 32'hFFFFFFF1;
    // rom_array[36886] = 32'hFFFFFFF1;
    // rom_array[36887] = 32'hFFFFFFF1;
    // rom_array[36888] = 32'hFFFFFFF1;
    // rom_array[36889] = 32'hFFFFFFF0;
    // rom_array[36890] = 32'hFFFFFFF0;
    // rom_array[36891] = 32'hFFFFFFF1;
    // rom_array[36892] = 32'hFFFFFFF1;
    // rom_array[36893] = 32'hFFFFFFF0;
    // rom_array[36894] = 32'hFFFFFFF0;
    // rom_array[36895] = 32'hFFFFFFF1;
    // rom_array[36896] = 32'hFFFFFFF1;
    // rom_array[36897] = 32'hFFFFFFF0;
    // rom_array[36898] = 32'hFFFFFFF0;
    // rom_array[36899] = 32'hFFFFFFF1;
    // rom_array[36900] = 32'hFFFFFFF1;
    // rom_array[36901] = 32'hFFFFFFF0;
    // rom_array[36902] = 32'hFFFFFFF0;
    // rom_array[36903] = 32'hFFFFFFF1;
    // rom_array[36904] = 32'hFFFFFFF1;
    // rom_array[36905] = 32'hFFFFFFF0;
    // rom_array[36906] = 32'hFFFFFFF0;
    // rom_array[36907] = 32'hFFFFFFF1;
    // rom_array[36908] = 32'hFFFFFFF1;
    // rom_array[36909] = 32'hFFFFFFF0;
    // rom_array[36910] = 32'hFFFFFFF0;
    // rom_array[36911] = 32'hFFFFFFF1;
    // rom_array[36912] = 32'hFFFFFFF1;
    // rom_array[36913] = 32'hFFFFFFF0;
    // rom_array[36914] = 32'hFFFFFFF0;
    // rom_array[36915] = 32'hFFFFFFF1;
    // rom_array[36916] = 32'hFFFFFFF1;
    // rom_array[36917] = 32'hFFFFFFF0;
    // rom_array[36918] = 32'hFFFFFFF0;
    // rom_array[36919] = 32'hFFFFFFF1;
    // rom_array[36920] = 32'hFFFFFFF1;
    // rom_array[36921] = 32'hFFFFFFF1;
    // rom_array[36922] = 32'hFFFFFFF1;
    // rom_array[36923] = 32'hFFFFFFF1;
    // rom_array[36924] = 32'hFFFFFFF1;
    // rom_array[36925] = 32'hFFFFFFF1;
    // rom_array[36926] = 32'hFFFFFFF1;
    // rom_array[36927] = 32'hFFFFFFF1;
    // rom_array[36928] = 32'hFFFFFFF1;
    // rom_array[36929] = 32'hFFFFFFF1;
    // rom_array[36930] = 32'hFFFFFFF1;
    // rom_array[36931] = 32'hFFFFFFF1;
    // rom_array[36932] = 32'hFFFFFFF1;
    // rom_array[36933] = 32'hFFFFFFF1;
    // rom_array[36934] = 32'hFFFFFFF1;
    // rom_array[36935] = 32'hFFFFFFF1;
    // rom_array[36936] = 32'hFFFFFFF1;
    // rom_array[36937] = 32'hFFFFFFF1;
    // rom_array[36938] = 32'hFFFFFFF1;
    // rom_array[36939] = 32'hFFFFFFF1;
    // rom_array[36940] = 32'hFFFFFFF1;
    // rom_array[36941] = 32'hFFFFFFF1;
    // rom_array[36942] = 32'hFFFFFFF1;
    // rom_array[36943] = 32'hFFFFFFF1;
    // rom_array[36944] = 32'hFFFFFFF1;
    // rom_array[36945] = 32'hFFFFFFF1;
    // rom_array[36946] = 32'hFFFFFFF1;
    // rom_array[36947] = 32'hFFFFFFF1;
    // rom_array[36948] = 32'hFFFFFFF1;
    // rom_array[36949] = 32'hFFFFFFF1;
    // rom_array[36950] = 32'hFFFFFFF1;
    // rom_array[36951] = 32'hFFFFFFF1;
    // rom_array[36952] = 32'hFFFFFFF1;
    // rom_array[36953] = 32'hFFFFFFF1;
    // rom_array[36954] = 32'hFFFFFFF1;
    // rom_array[36955] = 32'hFFFFFFF1;
    // rom_array[36956] = 32'hFFFFFFF1;
    // rom_array[36957] = 32'hFFFFFFF1;
    // rom_array[36958] = 32'hFFFFFFF1;
    // rom_array[36959] = 32'hFFFFFFF1;
    // rom_array[36960] = 32'hFFFFFFF1;
    // rom_array[36961] = 32'hFFFFFFF1;
    // rom_array[36962] = 32'hFFFFFFF1;
    // rom_array[36963] = 32'hFFFFFFF1;
    // rom_array[36964] = 32'hFFFFFFF1;
    // rom_array[36965] = 32'hFFFFFFF1;
    // rom_array[36966] = 32'hFFFFFFF1;
    // rom_array[36967] = 32'hFFFFFFF1;
    // rom_array[36968] = 32'hFFFFFFF1;
    // rom_array[36969] = 32'hFFFFFFF0;
    // rom_array[36970] = 32'hFFFFFFF0;
    // rom_array[36971] = 32'hFFFFFFF1;
    // rom_array[36972] = 32'hFFFFFFF1;
    // rom_array[36973] = 32'hFFFFFFF0;
    // rom_array[36974] = 32'hFFFFFFF0;
    // rom_array[36975] = 32'hFFFFFFF1;
    // rom_array[36976] = 32'hFFFFFFF1;
    // rom_array[36977] = 32'hFFFFFFF0;
    // rom_array[36978] = 32'hFFFFFFF0;
    // rom_array[36979] = 32'hFFFFFFF1;
    // rom_array[36980] = 32'hFFFFFFF1;
    // rom_array[36981] = 32'hFFFFFFF0;
    // rom_array[36982] = 32'hFFFFFFF0;
    // rom_array[36983] = 32'hFFFFFFF1;
    // rom_array[36984] = 32'hFFFFFFF1;
    // rom_array[36985] = 32'hFFFFFFF1;
    // rom_array[36986] = 32'hFFFFFFF1;
    // rom_array[36987] = 32'hFFFFFFF1;
    // rom_array[36988] = 32'hFFFFFFF1;
    // rom_array[36989] = 32'hFFFFFFF1;
    // rom_array[36990] = 32'hFFFFFFF1;
    // rom_array[36991] = 32'hFFFFFFF1;
    // rom_array[36992] = 32'hFFFFFFF1;
    // rom_array[36993] = 32'hFFFFFFF1;
    // rom_array[36994] = 32'hFFFFFFF1;
    // rom_array[36995] = 32'hFFFFFFF1;
    // rom_array[36996] = 32'hFFFFFFF1;
    // rom_array[36997] = 32'hFFFFFFF1;
    // rom_array[36998] = 32'hFFFFFFF1;
    // rom_array[36999] = 32'hFFFFFFF1;
    // rom_array[37000] = 32'hFFFFFFF1;
    // rom_array[37001] = 32'hFFFFFFF0;
    // rom_array[37002] = 32'hFFFFFFF0;
    // rom_array[37003] = 32'hFFFFFFF1;
    // rom_array[37004] = 32'hFFFFFFF1;
    // rom_array[37005] = 32'hFFFFFFF0;
    // rom_array[37006] = 32'hFFFFFFF0;
    // rom_array[37007] = 32'hFFFFFFF1;
    // rom_array[37008] = 32'hFFFFFFF1;
    // rom_array[37009] = 32'hFFFFFFF0;
    // rom_array[37010] = 32'hFFFFFFF0;
    // rom_array[37011] = 32'hFFFFFFF1;
    // rom_array[37012] = 32'hFFFFFFF1;
    // rom_array[37013] = 32'hFFFFFFF0;
    // rom_array[37014] = 32'hFFFFFFF0;
    // rom_array[37015] = 32'hFFFFFFF1;
    // rom_array[37016] = 32'hFFFFFFF1;
    // rom_array[37017] = 32'hFFFFFFF1;
    // rom_array[37018] = 32'hFFFFFFF1;
    // rom_array[37019] = 32'hFFFFFFF1;
    // rom_array[37020] = 32'hFFFFFFF1;
    // rom_array[37021] = 32'hFFFFFFF1;
    // rom_array[37022] = 32'hFFFFFFF1;
    // rom_array[37023] = 32'hFFFFFFF1;
    // rom_array[37024] = 32'hFFFFFFF1;
    // rom_array[37025] = 32'hFFFFFFF1;
    // rom_array[37026] = 32'hFFFFFFF1;
    // rom_array[37027] = 32'hFFFFFFF1;
    // rom_array[37028] = 32'hFFFFFFF1;
    // rom_array[37029] = 32'hFFFFFFF1;
    // rom_array[37030] = 32'hFFFFFFF1;
    // rom_array[37031] = 32'hFFFFFFF1;
    // rom_array[37032] = 32'hFFFFFFF1;
    // rom_array[37033] = 32'hFFFFFFF0;
    // rom_array[37034] = 32'hFFFFFFF0;
    // rom_array[37035] = 32'hFFFFFFF1;
    // rom_array[37036] = 32'hFFFFFFF1;
    // rom_array[37037] = 32'hFFFFFFF0;
    // rom_array[37038] = 32'hFFFFFFF0;
    // rom_array[37039] = 32'hFFFFFFF1;
    // rom_array[37040] = 32'hFFFFFFF1;
    // rom_array[37041] = 32'hFFFFFFF0;
    // rom_array[37042] = 32'hFFFFFFF0;
    // rom_array[37043] = 32'hFFFFFFF1;
    // rom_array[37044] = 32'hFFFFFFF1;
    // rom_array[37045] = 32'hFFFFFFF0;
    // rom_array[37046] = 32'hFFFFFFF0;
    // rom_array[37047] = 32'hFFFFFFF1;
    // rom_array[37048] = 32'hFFFFFFF1;
    // rom_array[37049] = 32'hFFFFFFF0;
    // rom_array[37050] = 32'hFFFFFFF0;
    // rom_array[37051] = 32'hFFFFFFF1;
    // rom_array[37052] = 32'hFFFFFFF1;
    // rom_array[37053] = 32'hFFFFFFF0;
    // rom_array[37054] = 32'hFFFFFFF0;
    // rom_array[37055] = 32'hFFFFFFF1;
    // rom_array[37056] = 32'hFFFFFFF1;
    // rom_array[37057] = 32'hFFFFFFF0;
    // rom_array[37058] = 32'hFFFFFFF0;
    // rom_array[37059] = 32'hFFFFFFF1;
    // rom_array[37060] = 32'hFFFFFFF1;
    // rom_array[37061] = 32'hFFFFFFF0;
    // rom_array[37062] = 32'hFFFFFFF0;
    // rom_array[37063] = 32'hFFFFFFF1;
    // rom_array[37064] = 32'hFFFFFFF1;
    // rom_array[37065] = 32'hFFFFFFF0;
    // rom_array[37066] = 32'hFFFFFFF0;
    // rom_array[37067] = 32'hFFFFFFF0;
    // rom_array[37068] = 32'hFFFFFFF0;
    // rom_array[37069] = 32'hFFFFFFF1;
    // rom_array[37070] = 32'hFFFFFFF1;
    // rom_array[37071] = 32'hFFFFFFF1;
    // rom_array[37072] = 32'hFFFFFFF1;
    // rom_array[37073] = 32'hFFFFFFF0;
    // rom_array[37074] = 32'hFFFFFFF0;
    // rom_array[37075] = 32'hFFFFFFF0;
    // rom_array[37076] = 32'hFFFFFFF0;
    // rom_array[37077] = 32'hFFFFFFF1;
    // rom_array[37078] = 32'hFFFFFFF1;
    // rom_array[37079] = 32'hFFFFFFF1;
    // rom_array[37080] = 32'hFFFFFFF1;
    // rom_array[37081] = 32'hFFFFFFF0;
    // rom_array[37082] = 32'hFFFFFFF0;
    // rom_array[37083] = 32'hFFFFFFF0;
    // rom_array[37084] = 32'hFFFFFFF0;
    // rom_array[37085] = 32'hFFFFFFF1;
    // rom_array[37086] = 32'hFFFFFFF1;
    // rom_array[37087] = 32'hFFFFFFF1;
    // rom_array[37088] = 32'hFFFFFFF1;
    // rom_array[37089] = 32'hFFFFFFF0;
    // rom_array[37090] = 32'hFFFFFFF0;
    // rom_array[37091] = 32'hFFFFFFF0;
    // rom_array[37092] = 32'hFFFFFFF0;
    // rom_array[37093] = 32'hFFFFFFF1;
    // rom_array[37094] = 32'hFFFFFFF1;
    // rom_array[37095] = 32'hFFFFFFF1;
    // rom_array[37096] = 32'hFFFFFFF1;
    // rom_array[37097] = 32'hFFFFFFF0;
    // rom_array[37098] = 32'hFFFFFFF0;
    // rom_array[37099] = 32'hFFFFFFF0;
    // rom_array[37100] = 32'hFFFFFFF0;
    // rom_array[37101] = 32'hFFFFFFF1;
    // rom_array[37102] = 32'hFFFFFFF1;
    // rom_array[37103] = 32'hFFFFFFF1;
    // rom_array[37104] = 32'hFFFFFFF1;
    // rom_array[37105] = 32'hFFFFFFF0;
    // rom_array[37106] = 32'hFFFFFFF0;
    // rom_array[37107] = 32'hFFFFFFF0;
    // rom_array[37108] = 32'hFFFFFFF0;
    // rom_array[37109] = 32'hFFFFFFF1;
    // rom_array[37110] = 32'hFFFFFFF1;
    // rom_array[37111] = 32'hFFFFFFF1;
    // rom_array[37112] = 32'hFFFFFFF1;
    // rom_array[37113] = 32'hFFFFFFF0;
    // rom_array[37114] = 32'hFFFFFFF0;
    // rom_array[37115] = 32'hFFFFFFF0;
    // rom_array[37116] = 32'hFFFFFFF0;
    // rom_array[37117] = 32'hFFFFFFF1;
    // rom_array[37118] = 32'hFFFFFFF1;
    // rom_array[37119] = 32'hFFFFFFF1;
    // rom_array[37120] = 32'hFFFFFFF1;
    // rom_array[37121] = 32'hFFFFFFF0;
    // rom_array[37122] = 32'hFFFFFFF0;
    // rom_array[37123] = 32'hFFFFFFF0;
    // rom_array[37124] = 32'hFFFFFFF0;
    // rom_array[37125] = 32'hFFFFFFF1;
    // rom_array[37126] = 32'hFFFFFFF1;
    // rom_array[37127] = 32'hFFFFFFF1;
    // rom_array[37128] = 32'hFFFFFFF1;
    // rom_array[37129] = 32'hFFFFFFF0;
    // rom_array[37130] = 32'hFFFFFFF0;
    // rom_array[37131] = 32'hFFFFFFF0;
    // rom_array[37132] = 32'hFFFFFFF0;
    // rom_array[37133] = 32'hFFFFFFF1;
    // rom_array[37134] = 32'hFFFFFFF1;
    // rom_array[37135] = 32'hFFFFFFF1;
    // rom_array[37136] = 32'hFFFFFFF1;
    // rom_array[37137] = 32'hFFFFFFF0;
    // rom_array[37138] = 32'hFFFFFFF0;
    // rom_array[37139] = 32'hFFFFFFF0;
    // rom_array[37140] = 32'hFFFFFFF0;
    // rom_array[37141] = 32'hFFFFFFF1;
    // rom_array[37142] = 32'hFFFFFFF1;
    // rom_array[37143] = 32'hFFFFFFF1;
    // rom_array[37144] = 32'hFFFFFFF1;
    // rom_array[37145] = 32'hFFFFFFF0;
    // rom_array[37146] = 32'hFFFFFFF0;
    // rom_array[37147] = 32'hFFFFFFF0;
    // rom_array[37148] = 32'hFFFFFFF0;
    // rom_array[37149] = 32'hFFFFFFF1;
    // rom_array[37150] = 32'hFFFFFFF1;
    // rom_array[37151] = 32'hFFFFFFF1;
    // rom_array[37152] = 32'hFFFFFFF1;
    // rom_array[37153] = 32'hFFFFFFF0;
    // rom_array[37154] = 32'hFFFFFFF0;
    // rom_array[37155] = 32'hFFFFFFF0;
    // rom_array[37156] = 32'hFFFFFFF0;
    // rom_array[37157] = 32'hFFFFFFF1;
    // rom_array[37158] = 32'hFFFFFFF1;
    // rom_array[37159] = 32'hFFFFFFF1;
    // rom_array[37160] = 32'hFFFFFFF1;
    // rom_array[37161] = 32'hFFFFFFF0;
    // rom_array[37162] = 32'hFFFFFFF0;
    // rom_array[37163] = 32'hFFFFFFF0;
    // rom_array[37164] = 32'hFFFFFFF0;
    // rom_array[37165] = 32'hFFFFFFF1;
    // rom_array[37166] = 32'hFFFFFFF1;
    // rom_array[37167] = 32'hFFFFFFF1;
    // rom_array[37168] = 32'hFFFFFFF1;
    // rom_array[37169] = 32'hFFFFFFF0;
    // rom_array[37170] = 32'hFFFFFFF0;
    // rom_array[37171] = 32'hFFFFFFF0;
    // rom_array[37172] = 32'hFFFFFFF0;
    // rom_array[37173] = 32'hFFFFFFF1;
    // rom_array[37174] = 32'hFFFFFFF1;
    // rom_array[37175] = 32'hFFFFFFF1;
    // rom_array[37176] = 32'hFFFFFFF1;
    // rom_array[37177] = 32'hFFFFFFF0;
    // rom_array[37178] = 32'hFFFFFFF0;
    // rom_array[37179] = 32'hFFFFFFF0;
    // rom_array[37180] = 32'hFFFFFFF0;
    // rom_array[37181] = 32'hFFFFFFF1;
    // rom_array[37182] = 32'hFFFFFFF1;
    // rom_array[37183] = 32'hFFFFFFF1;
    // rom_array[37184] = 32'hFFFFFFF1;
    // rom_array[37185] = 32'hFFFFFFF0;
    // rom_array[37186] = 32'hFFFFFFF0;
    // rom_array[37187] = 32'hFFFFFFF0;
    // rom_array[37188] = 32'hFFFFFFF0;
    // rom_array[37189] = 32'hFFFFFFF1;
    // rom_array[37190] = 32'hFFFFFFF1;
    // rom_array[37191] = 32'hFFFFFFF1;
    // rom_array[37192] = 32'hFFFFFFF1;
    // rom_array[37193] = 32'hFFFFFFF0;
    // rom_array[37194] = 32'hFFFFFFF0;
    // rom_array[37195] = 32'hFFFFFFF0;
    // rom_array[37196] = 32'hFFFFFFF0;
    // rom_array[37197] = 32'hFFFFFFF0;
    // rom_array[37198] = 32'hFFFFFFF0;
    // rom_array[37199] = 32'hFFFFFFF1;
    // rom_array[37200] = 32'hFFFFFFF1;
    // rom_array[37201] = 32'hFFFFFFF0;
    // rom_array[37202] = 32'hFFFFFFF0;
    // rom_array[37203] = 32'hFFFFFFF0;
    // rom_array[37204] = 32'hFFFFFFF0;
    // rom_array[37205] = 32'hFFFFFFF0;
    // rom_array[37206] = 32'hFFFFFFF0;
    // rom_array[37207] = 32'hFFFFFFF1;
    // rom_array[37208] = 32'hFFFFFFF1;
    // rom_array[37209] = 32'hFFFFFFF0;
    // rom_array[37210] = 32'hFFFFFFF0;
    // rom_array[37211] = 32'hFFFFFFF0;
    // rom_array[37212] = 32'hFFFFFFF0;
    // rom_array[37213] = 32'hFFFFFFF1;
    // rom_array[37214] = 32'hFFFFFFF1;
    // rom_array[37215] = 32'hFFFFFFF1;
    // rom_array[37216] = 32'hFFFFFFF1;
    // rom_array[37217] = 32'hFFFFFFF0;
    // rom_array[37218] = 32'hFFFFFFF0;
    // rom_array[37219] = 32'hFFFFFFF0;
    // rom_array[37220] = 32'hFFFFFFF0;
    // rom_array[37221] = 32'hFFFFFFF1;
    // rom_array[37222] = 32'hFFFFFFF1;
    // rom_array[37223] = 32'hFFFFFFF1;
    // rom_array[37224] = 32'hFFFFFFF1;
    // rom_array[37225] = 32'hFFFFFFF0;
    // rom_array[37226] = 32'hFFFFFFF0;
    // rom_array[37227] = 32'hFFFFFFF0;
    // rom_array[37228] = 32'hFFFFFFF0;
    // rom_array[37229] = 32'hFFFFFFF1;
    // rom_array[37230] = 32'hFFFFFFF1;
    // rom_array[37231] = 32'hFFFFFFF1;
    // rom_array[37232] = 32'hFFFFFFF1;
    // rom_array[37233] = 32'hFFFFFFF0;
    // rom_array[37234] = 32'hFFFFFFF0;
    // rom_array[37235] = 32'hFFFFFFF0;
    // rom_array[37236] = 32'hFFFFFFF0;
    // rom_array[37237] = 32'hFFFFFFF1;
    // rom_array[37238] = 32'hFFFFFFF1;
    // rom_array[37239] = 32'hFFFFFFF1;
    // rom_array[37240] = 32'hFFFFFFF1;
    // rom_array[37241] = 32'hFFFFFFF0;
    // rom_array[37242] = 32'hFFFFFFF0;
    // rom_array[37243] = 32'hFFFFFFF0;
    // rom_array[37244] = 32'hFFFFFFF0;
    // rom_array[37245] = 32'hFFFFFFF1;
    // rom_array[37246] = 32'hFFFFFFF1;
    // rom_array[37247] = 32'hFFFFFFF1;
    // rom_array[37248] = 32'hFFFFFFF1;
    // rom_array[37249] = 32'hFFFFFFF0;
    // rom_array[37250] = 32'hFFFFFFF0;
    // rom_array[37251] = 32'hFFFFFFF0;
    // rom_array[37252] = 32'hFFFFFFF0;
    // rom_array[37253] = 32'hFFFFFFF1;
    // rom_array[37254] = 32'hFFFFFFF1;
    // rom_array[37255] = 32'hFFFFFFF1;
    // rom_array[37256] = 32'hFFFFFFF1;
    // rom_array[37257] = 32'hFFFFFFF0;
    // rom_array[37258] = 32'hFFFFFFF0;
    // rom_array[37259] = 32'hFFFFFFF1;
    // rom_array[37260] = 32'hFFFFFFF1;
    // rom_array[37261] = 32'hFFFFFFF0;
    // rom_array[37262] = 32'hFFFFFFF0;
    // rom_array[37263] = 32'hFFFFFFF1;
    // rom_array[37264] = 32'hFFFFFFF1;
    // rom_array[37265] = 32'hFFFFFFF0;
    // rom_array[37266] = 32'hFFFFFFF0;
    // rom_array[37267] = 32'hFFFFFFF1;
    // rom_array[37268] = 32'hFFFFFFF1;
    // rom_array[37269] = 32'hFFFFFFF0;
    // rom_array[37270] = 32'hFFFFFFF0;
    // rom_array[37271] = 32'hFFFFFFF1;
    // rom_array[37272] = 32'hFFFFFFF1;
    // rom_array[37273] = 32'hFFFFFFF0;
    // rom_array[37274] = 32'hFFFFFFF0;
    // rom_array[37275] = 32'hFFFFFFF1;
    // rom_array[37276] = 32'hFFFFFFF1;
    // rom_array[37277] = 32'hFFFFFFF0;
    // rom_array[37278] = 32'hFFFFFFF0;
    // rom_array[37279] = 32'hFFFFFFF1;
    // rom_array[37280] = 32'hFFFFFFF1;
    // rom_array[37281] = 32'hFFFFFFF0;
    // rom_array[37282] = 32'hFFFFFFF0;
    // rom_array[37283] = 32'hFFFFFFF1;
    // rom_array[37284] = 32'hFFFFFFF1;
    // rom_array[37285] = 32'hFFFFFFF0;
    // rom_array[37286] = 32'hFFFFFFF0;
    // rom_array[37287] = 32'hFFFFFFF1;
    // rom_array[37288] = 32'hFFFFFFF1;
    // rom_array[37289] = 32'hFFFFFFF0;
    // rom_array[37290] = 32'hFFFFFFF0;
    // rom_array[37291] = 32'hFFFFFFF0;
    // rom_array[37292] = 32'hFFFFFFF0;
    // rom_array[37293] = 32'hFFFFFFF1;
    // rom_array[37294] = 32'hFFFFFFF1;
    // rom_array[37295] = 32'hFFFFFFF1;
    // rom_array[37296] = 32'hFFFFFFF1;
    // rom_array[37297] = 32'hFFFFFFF0;
    // rom_array[37298] = 32'hFFFFFFF0;
    // rom_array[37299] = 32'hFFFFFFF0;
    // rom_array[37300] = 32'hFFFFFFF0;
    // rom_array[37301] = 32'hFFFFFFF1;
    // rom_array[37302] = 32'hFFFFFFF1;
    // rom_array[37303] = 32'hFFFFFFF1;
    // rom_array[37304] = 32'hFFFFFFF1;
    // rom_array[37305] = 32'hFFFFFFF1;
    // rom_array[37306] = 32'hFFFFFFF1;
    // rom_array[37307] = 32'hFFFFFFF1;
    // rom_array[37308] = 32'hFFFFFFF1;
    // rom_array[37309] = 32'hFFFFFFF1;
    // rom_array[37310] = 32'hFFFFFFF1;
    // rom_array[37311] = 32'hFFFFFFF1;
    // rom_array[37312] = 32'hFFFFFFF1;
    // rom_array[37313] = 32'hFFFFFFF1;
    // rom_array[37314] = 32'hFFFFFFF1;
    // rom_array[37315] = 32'hFFFFFFF1;
    // rom_array[37316] = 32'hFFFFFFF1;
    // rom_array[37317] = 32'hFFFFFFF1;
    // rom_array[37318] = 32'hFFFFFFF1;
    // rom_array[37319] = 32'hFFFFFFF1;
    // rom_array[37320] = 32'hFFFFFFF1;
    // rom_array[37321] = 32'hFFFFFFF1;
    // rom_array[37322] = 32'hFFFFFFF1;
    // rom_array[37323] = 32'hFFFFFFF1;
    // rom_array[37324] = 32'hFFFFFFF1;
    // rom_array[37325] = 32'hFFFFFFF1;
    // rom_array[37326] = 32'hFFFFFFF1;
    // rom_array[37327] = 32'hFFFFFFF1;
    // rom_array[37328] = 32'hFFFFFFF1;
    // rom_array[37329] = 32'hFFFFFFF1;
    // rom_array[37330] = 32'hFFFFFFF1;
    // rom_array[37331] = 32'hFFFFFFF1;
    // rom_array[37332] = 32'hFFFFFFF1;
    // rom_array[37333] = 32'hFFFFFFF1;
    // rom_array[37334] = 32'hFFFFFFF1;
    // rom_array[37335] = 32'hFFFFFFF1;
    // rom_array[37336] = 32'hFFFFFFF1;
    // rom_array[37337] = 32'hFFFFFFF0;
    // rom_array[37338] = 32'hFFFFFFF0;
    // rom_array[37339] = 32'hFFFFFFF1;
    // rom_array[37340] = 32'hFFFFFFF1;
    // rom_array[37341] = 32'hFFFFFFF0;
    // rom_array[37342] = 32'hFFFFFFF0;
    // rom_array[37343] = 32'hFFFFFFF1;
    // rom_array[37344] = 32'hFFFFFFF1;
    // rom_array[37345] = 32'hFFFFFFF0;
    // rom_array[37346] = 32'hFFFFFFF0;
    // rom_array[37347] = 32'hFFFFFFF1;
    // rom_array[37348] = 32'hFFFFFFF1;
    // rom_array[37349] = 32'hFFFFFFF0;
    // rom_array[37350] = 32'hFFFFFFF0;
    // rom_array[37351] = 32'hFFFFFFF1;
    // rom_array[37352] = 32'hFFFFFFF1;
    // rom_array[37353] = 32'hFFFFFFF0;
    // rom_array[37354] = 32'hFFFFFFF0;
    // rom_array[37355] = 32'hFFFFFFF0;
    // rom_array[37356] = 32'hFFFFFFF0;
    // rom_array[37357] = 32'hFFFFFFF1;
    // rom_array[37358] = 32'hFFFFFFF1;
    // rom_array[37359] = 32'hFFFFFFF1;
    // rom_array[37360] = 32'hFFFFFFF1;
    // rom_array[37361] = 32'hFFFFFFF0;
    // rom_array[37362] = 32'hFFFFFFF0;
    // rom_array[37363] = 32'hFFFFFFF0;
    // rom_array[37364] = 32'hFFFFFFF0;
    // rom_array[37365] = 32'hFFFFFFF1;
    // rom_array[37366] = 32'hFFFFFFF1;
    // rom_array[37367] = 32'hFFFFFFF1;
    // rom_array[37368] = 32'hFFFFFFF1;
    // rom_array[37369] = 32'hFFFFFFF0;
    // rom_array[37370] = 32'hFFFFFFF0;
    // rom_array[37371] = 32'hFFFFFFF1;
    // rom_array[37372] = 32'hFFFFFFF1;
    // rom_array[37373] = 32'hFFFFFFF0;
    // rom_array[37374] = 32'hFFFFFFF0;
    // rom_array[37375] = 32'hFFFFFFF1;
    // rom_array[37376] = 32'hFFFFFFF1;
    // rom_array[37377] = 32'hFFFFFFF0;
    // rom_array[37378] = 32'hFFFFFFF0;
    // rom_array[37379] = 32'hFFFFFFF1;
    // rom_array[37380] = 32'hFFFFFFF1;
    // rom_array[37381] = 32'hFFFFFFF0;
    // rom_array[37382] = 32'hFFFFFFF0;
    // rom_array[37383] = 32'hFFFFFFF1;
    // rom_array[37384] = 32'hFFFFFFF1;
    // rom_array[37385] = 32'hFFFFFFF0;
    // rom_array[37386] = 32'hFFFFFFF0;
    // rom_array[37387] = 32'hFFFFFFF0;
    // rom_array[37388] = 32'hFFFFFFF0;
    // rom_array[37389] = 32'hFFFFFFF1;
    // rom_array[37390] = 32'hFFFFFFF1;
    // rom_array[37391] = 32'hFFFFFFF1;
    // rom_array[37392] = 32'hFFFFFFF1;
    // rom_array[37393] = 32'hFFFFFFF0;
    // rom_array[37394] = 32'hFFFFFFF0;
    // rom_array[37395] = 32'hFFFFFFF0;
    // rom_array[37396] = 32'hFFFFFFF0;
    // rom_array[37397] = 32'hFFFFFFF1;
    // rom_array[37398] = 32'hFFFFFFF1;
    // rom_array[37399] = 32'hFFFFFFF1;
    // rom_array[37400] = 32'hFFFFFFF1;
    // rom_array[37401] = 32'hFFFFFFF0;
    // rom_array[37402] = 32'hFFFFFFF0;
    // rom_array[37403] = 32'hFFFFFFF0;
    // rom_array[37404] = 32'hFFFFFFF0;
    // rom_array[37405] = 32'hFFFFFFF1;
    // rom_array[37406] = 32'hFFFFFFF1;
    // rom_array[37407] = 32'hFFFFFFF1;
    // rom_array[37408] = 32'hFFFFFFF1;
    // rom_array[37409] = 32'hFFFFFFF0;
    // rom_array[37410] = 32'hFFFFFFF0;
    // rom_array[37411] = 32'hFFFFFFF0;
    // rom_array[37412] = 32'hFFFFFFF0;
    // rom_array[37413] = 32'hFFFFFFF1;
    // rom_array[37414] = 32'hFFFFFFF1;
    // rom_array[37415] = 32'hFFFFFFF1;
    // rom_array[37416] = 32'hFFFFFFF1;
    // rom_array[37417] = 32'hFFFFFFF0;
    // rom_array[37418] = 32'hFFFFFFF0;
    // rom_array[37419] = 32'hFFFFFFF1;
    // rom_array[37420] = 32'hFFFFFFF1;
    // rom_array[37421] = 32'hFFFFFFF0;
    // rom_array[37422] = 32'hFFFFFFF0;
    // rom_array[37423] = 32'hFFFFFFF1;
    // rom_array[37424] = 32'hFFFFFFF1;
    // rom_array[37425] = 32'hFFFFFFF0;
    // rom_array[37426] = 32'hFFFFFFF0;
    // rom_array[37427] = 32'hFFFFFFF1;
    // rom_array[37428] = 32'hFFFFFFF1;
    // rom_array[37429] = 32'hFFFFFFF0;
    // rom_array[37430] = 32'hFFFFFFF0;
    // rom_array[37431] = 32'hFFFFFFF1;
    // rom_array[37432] = 32'hFFFFFFF1;
    // rom_array[37433] = 32'hFFFFFFF0;
    // rom_array[37434] = 32'hFFFFFFF0;
    // rom_array[37435] = 32'hFFFFFFF1;
    // rom_array[37436] = 32'hFFFFFFF1;
    // rom_array[37437] = 32'hFFFFFFF0;
    // rom_array[37438] = 32'hFFFFFFF0;
    // rom_array[37439] = 32'hFFFFFFF1;
    // rom_array[37440] = 32'hFFFFFFF1;
    // rom_array[37441] = 32'hFFFFFFF0;
    // rom_array[37442] = 32'hFFFFFFF0;
    // rom_array[37443] = 32'hFFFFFFF1;
    // rom_array[37444] = 32'hFFFFFFF1;
    // rom_array[37445] = 32'hFFFFFFF0;
    // rom_array[37446] = 32'hFFFFFFF0;
    // rom_array[37447] = 32'hFFFFFFF1;
    // rom_array[37448] = 32'hFFFFFFF1;
    // rom_array[37449] = 32'hFFFFFFF0;
    // rom_array[37450] = 32'hFFFFFFF0;
    // rom_array[37451] = 32'hFFFFFFF1;
    // rom_array[37452] = 32'hFFFFFFF1;
    // rom_array[37453] = 32'hFFFFFFF0;
    // rom_array[37454] = 32'hFFFFFFF0;
    // rom_array[37455] = 32'hFFFFFFF1;
    // rom_array[37456] = 32'hFFFFFFF1;
    // rom_array[37457] = 32'hFFFFFFF0;
    // rom_array[37458] = 32'hFFFFFFF0;
    // rom_array[37459] = 32'hFFFFFFF1;
    // rom_array[37460] = 32'hFFFFFFF1;
    // rom_array[37461] = 32'hFFFFFFF0;
    // rom_array[37462] = 32'hFFFFFFF0;
    // rom_array[37463] = 32'hFFFFFFF1;
    // rom_array[37464] = 32'hFFFFFFF1;
    // rom_array[37465] = 32'hFFFFFFF1;
    // rom_array[37466] = 32'hFFFFFFF1;
    // rom_array[37467] = 32'hFFFFFFF1;
    // rom_array[37468] = 32'hFFFFFFF1;
    // rom_array[37469] = 32'hFFFFFFF0;
    // rom_array[37470] = 32'hFFFFFFF0;
    // rom_array[37471] = 32'hFFFFFFF0;
    // rom_array[37472] = 32'hFFFFFFF0;
    // rom_array[37473] = 32'hFFFFFFF1;
    // rom_array[37474] = 32'hFFFFFFF1;
    // rom_array[37475] = 32'hFFFFFFF1;
    // rom_array[37476] = 32'hFFFFFFF1;
    // rom_array[37477] = 32'hFFFFFFF0;
    // rom_array[37478] = 32'hFFFFFFF0;
    // rom_array[37479] = 32'hFFFFFFF0;
    // rom_array[37480] = 32'hFFFFFFF0;
    // rom_array[37481] = 32'hFFFFFFF0;
    // rom_array[37482] = 32'hFFFFFFF0;
    // rom_array[37483] = 32'hFFFFFFF1;
    // rom_array[37484] = 32'hFFFFFFF1;
    // rom_array[37485] = 32'hFFFFFFF0;
    // rom_array[37486] = 32'hFFFFFFF0;
    // rom_array[37487] = 32'hFFFFFFF1;
    // rom_array[37488] = 32'hFFFFFFF1;
    // rom_array[37489] = 32'hFFFFFFF0;
    // rom_array[37490] = 32'hFFFFFFF0;
    // rom_array[37491] = 32'hFFFFFFF1;
    // rom_array[37492] = 32'hFFFFFFF1;
    // rom_array[37493] = 32'hFFFFFFF0;
    // rom_array[37494] = 32'hFFFFFFF0;
    // rom_array[37495] = 32'hFFFFFFF1;
    // rom_array[37496] = 32'hFFFFFFF1;
    // rom_array[37497] = 32'hFFFFFFF1;
    // rom_array[37498] = 32'hFFFFFFF1;
    // rom_array[37499] = 32'hFFFFFFF1;
    // rom_array[37500] = 32'hFFFFFFF1;
    // rom_array[37501] = 32'hFFFFFFF0;
    // rom_array[37502] = 32'hFFFFFFF0;
    // rom_array[37503] = 32'hFFFFFFF0;
    // rom_array[37504] = 32'hFFFFFFF0;
    // rom_array[37505] = 32'hFFFFFFF1;
    // rom_array[37506] = 32'hFFFFFFF1;
    // rom_array[37507] = 32'hFFFFFFF1;
    // rom_array[37508] = 32'hFFFFFFF1;
    // rom_array[37509] = 32'hFFFFFFF0;
    // rom_array[37510] = 32'hFFFFFFF0;
    // rom_array[37511] = 32'hFFFFFFF0;
    // rom_array[37512] = 32'hFFFFFFF0;
    // rom_array[37513] = 32'hFFFFFFF1;
    // rom_array[37514] = 32'hFFFFFFF1;
    // rom_array[37515] = 32'hFFFFFFF1;
    // rom_array[37516] = 32'hFFFFFFF1;
    // rom_array[37517] = 32'hFFFFFFF0;
    // rom_array[37518] = 32'hFFFFFFF0;
    // rom_array[37519] = 32'hFFFFFFF0;
    // rom_array[37520] = 32'hFFFFFFF0;
    // rom_array[37521] = 32'hFFFFFFF1;
    // rom_array[37522] = 32'hFFFFFFF1;
    // rom_array[37523] = 32'hFFFFFFF1;
    // rom_array[37524] = 32'hFFFFFFF1;
    // rom_array[37525] = 32'hFFFFFFF0;
    // rom_array[37526] = 32'hFFFFFFF0;
    // rom_array[37527] = 32'hFFFFFFF0;
    // rom_array[37528] = 32'hFFFFFFF0;
    // rom_array[37529] = 32'hFFFFFFF0;
    // rom_array[37530] = 32'hFFFFFFF0;
    // rom_array[37531] = 32'hFFFFFFF1;
    // rom_array[37532] = 32'hFFFFFFF1;
    // rom_array[37533] = 32'hFFFFFFF0;
    // rom_array[37534] = 32'hFFFFFFF0;
    // rom_array[37535] = 32'hFFFFFFF1;
    // rom_array[37536] = 32'hFFFFFFF1;
    // rom_array[37537] = 32'hFFFFFFF0;
    // rom_array[37538] = 32'hFFFFFFF0;
    // rom_array[37539] = 32'hFFFFFFF1;
    // rom_array[37540] = 32'hFFFFFFF1;
    // rom_array[37541] = 32'hFFFFFFF0;
    // rom_array[37542] = 32'hFFFFFFF0;
    // rom_array[37543] = 32'hFFFFFFF1;
    // rom_array[37544] = 32'hFFFFFFF1;
    // rom_array[37545] = 32'hFFFFFFF0;
    // rom_array[37546] = 32'hFFFFFFF0;
    // rom_array[37547] = 32'hFFFFFFF1;
    // rom_array[37548] = 32'hFFFFFFF1;
    // rom_array[37549] = 32'hFFFFFFF0;
    // rom_array[37550] = 32'hFFFFFFF0;
    // rom_array[37551] = 32'hFFFFFFF1;
    // rom_array[37552] = 32'hFFFFFFF1;
    // rom_array[37553] = 32'hFFFFFFF0;
    // rom_array[37554] = 32'hFFFFFFF0;
    // rom_array[37555] = 32'hFFFFFFF1;
    // rom_array[37556] = 32'hFFFFFFF1;
    // rom_array[37557] = 32'hFFFFFFF0;
    // rom_array[37558] = 32'hFFFFFFF0;
    // rom_array[37559] = 32'hFFFFFFF1;
    // rom_array[37560] = 32'hFFFFFFF1;
    // rom_array[37561] = 32'hFFFFFFF0;
    // rom_array[37562] = 32'hFFFFFFF0;
    // rom_array[37563] = 32'hFFFFFFF1;
    // rom_array[37564] = 32'hFFFFFFF1;
    // rom_array[37565] = 32'hFFFFFFF1;
    // rom_array[37566] = 32'hFFFFFFF1;
    // rom_array[37567] = 32'hFFFFFFF1;
    // rom_array[37568] = 32'hFFFFFFF1;
    // rom_array[37569] = 32'hFFFFFFF0;
    // rom_array[37570] = 32'hFFFFFFF0;
    // rom_array[37571] = 32'hFFFFFFF1;
    // rom_array[37572] = 32'hFFFFFFF1;
    // rom_array[37573] = 32'hFFFFFFF1;
    // rom_array[37574] = 32'hFFFFFFF1;
    // rom_array[37575] = 32'hFFFFFFF1;
    // rom_array[37576] = 32'hFFFFFFF1;
    // rom_array[37577] = 32'hFFFFFFF0;
    // rom_array[37578] = 32'hFFFFFFF0;
    // rom_array[37579] = 32'hFFFFFFF0;
    // rom_array[37580] = 32'hFFFFFFF0;
    // rom_array[37581] = 32'hFFFFFFF1;
    // rom_array[37582] = 32'hFFFFFFF1;
    // rom_array[37583] = 32'hFFFFFFF1;
    // rom_array[37584] = 32'hFFFFFFF1;
    // rom_array[37585] = 32'hFFFFFFF0;
    // rom_array[37586] = 32'hFFFFFFF0;
    // rom_array[37587] = 32'hFFFFFFF0;
    // rom_array[37588] = 32'hFFFFFFF0;
    // rom_array[37589] = 32'hFFFFFFF1;
    // rom_array[37590] = 32'hFFFFFFF1;
    // rom_array[37591] = 32'hFFFFFFF1;
    // rom_array[37592] = 32'hFFFFFFF1;
    // rom_array[37593] = 32'hFFFFFFF0;
    // rom_array[37594] = 32'hFFFFFFF0;
    // rom_array[37595] = 32'hFFFFFFF1;
    // rom_array[37596] = 32'hFFFFFFF1;
    // rom_array[37597] = 32'hFFFFFFF0;
    // rom_array[37598] = 32'hFFFFFFF0;
    // rom_array[37599] = 32'hFFFFFFF1;
    // rom_array[37600] = 32'hFFFFFFF1;
    // rom_array[37601] = 32'hFFFFFFF0;
    // rom_array[37602] = 32'hFFFFFFF0;
    // rom_array[37603] = 32'hFFFFFFF1;
    // rom_array[37604] = 32'hFFFFFFF1;
    // rom_array[37605] = 32'hFFFFFFF0;
    // rom_array[37606] = 32'hFFFFFFF0;
    // rom_array[37607] = 32'hFFFFFFF1;
    // rom_array[37608] = 32'hFFFFFFF1;
    // rom_array[37609] = 32'hFFFFFFF0;
    // rom_array[37610] = 32'hFFFFFFF0;
    // rom_array[37611] = 32'hFFFFFFF0;
    // rom_array[37612] = 32'hFFFFFFF0;
    // rom_array[37613] = 32'hFFFFFFF1;
    // rom_array[37614] = 32'hFFFFFFF1;
    // rom_array[37615] = 32'hFFFFFFF1;
    // rom_array[37616] = 32'hFFFFFFF1;
    // rom_array[37617] = 32'hFFFFFFF0;
    // rom_array[37618] = 32'hFFFFFFF0;
    // rom_array[37619] = 32'hFFFFFFF0;
    // rom_array[37620] = 32'hFFFFFFF0;
    // rom_array[37621] = 32'hFFFFFFF1;
    // rom_array[37622] = 32'hFFFFFFF1;
    // rom_array[37623] = 32'hFFFFFFF1;
    // rom_array[37624] = 32'hFFFFFFF1;
    // rom_array[37625] = 32'hFFFFFFF0;
    // rom_array[37626] = 32'hFFFFFFF0;
    // rom_array[37627] = 32'hFFFFFFF0;
    // rom_array[37628] = 32'hFFFFFFF0;
    // rom_array[37629] = 32'hFFFFFFF1;
    // rom_array[37630] = 32'hFFFFFFF1;
    // rom_array[37631] = 32'hFFFFFFF1;
    // rom_array[37632] = 32'hFFFFFFF1;
    // rom_array[37633] = 32'hFFFFFFF0;
    // rom_array[37634] = 32'hFFFFFFF0;
    // rom_array[37635] = 32'hFFFFFFF0;
    // rom_array[37636] = 32'hFFFFFFF0;
    // rom_array[37637] = 32'hFFFFFFF1;
    // rom_array[37638] = 32'hFFFFFFF1;
    // rom_array[37639] = 32'hFFFFFFF1;
    // rom_array[37640] = 32'hFFFFFFF1;
    // rom_array[37641] = 32'hFFFFFFF0;
    // rom_array[37642] = 32'hFFFFFFF0;
    // rom_array[37643] = 32'hFFFFFFF1;
    // rom_array[37644] = 32'hFFFFFFF1;
    // rom_array[37645] = 32'hFFFFFFF0;
    // rom_array[37646] = 32'hFFFFFFF0;
    // rom_array[37647] = 32'hFFFFFFF1;
    // rom_array[37648] = 32'hFFFFFFF1;
    // rom_array[37649] = 32'hFFFFFFF0;
    // rom_array[37650] = 32'hFFFFFFF0;
    // rom_array[37651] = 32'hFFFFFFF1;
    // rom_array[37652] = 32'hFFFFFFF1;
    // rom_array[37653] = 32'hFFFFFFF0;
    // rom_array[37654] = 32'hFFFFFFF0;
    // rom_array[37655] = 32'hFFFFFFF1;
    // rom_array[37656] = 32'hFFFFFFF1;
    // rom_array[37657] = 32'hFFFFFFF0;
    // rom_array[37658] = 32'hFFFFFFF0;
    // rom_array[37659] = 32'hFFFFFFF1;
    // rom_array[37660] = 32'hFFFFFFF1;
    // rom_array[37661] = 32'hFFFFFFF0;
    // rom_array[37662] = 32'hFFFFFFF0;
    // rom_array[37663] = 32'hFFFFFFF1;
    // rom_array[37664] = 32'hFFFFFFF1;
    // rom_array[37665] = 32'hFFFFFFF0;
    // rom_array[37666] = 32'hFFFFFFF0;
    // rom_array[37667] = 32'hFFFFFFF1;
    // rom_array[37668] = 32'hFFFFFFF1;
    // rom_array[37669] = 32'hFFFFFFF0;
    // rom_array[37670] = 32'hFFFFFFF0;
    // rom_array[37671] = 32'hFFFFFFF1;
    // rom_array[37672] = 32'hFFFFFFF1;
    // rom_array[37673] = 32'hFFFFFFF1;
    // rom_array[37674] = 32'hFFFFFFF1;
    // rom_array[37675] = 32'hFFFFFFF1;
    // rom_array[37676] = 32'hFFFFFFF1;
    // rom_array[37677] = 32'hFFFFFFF1;
    // rom_array[37678] = 32'hFFFFFFF1;
    // rom_array[37679] = 32'hFFFFFFF1;
    // rom_array[37680] = 32'hFFFFFFF1;
    // rom_array[37681] = 32'hFFFFFFF1;
    // rom_array[37682] = 32'hFFFFFFF1;
    // rom_array[37683] = 32'hFFFFFFF1;
    // rom_array[37684] = 32'hFFFFFFF1;
    // rom_array[37685] = 32'hFFFFFFF1;
    // rom_array[37686] = 32'hFFFFFFF1;
    // rom_array[37687] = 32'hFFFFFFF1;
    // rom_array[37688] = 32'hFFFFFFF1;
    // rom_array[37689] = 32'hFFFFFFF0;
    // rom_array[37690] = 32'hFFFFFFF0;
    // rom_array[37691] = 32'hFFFFFFF0;
    // rom_array[37692] = 32'hFFFFFFF0;
    // rom_array[37693] = 32'hFFFFFFF1;
    // rom_array[37694] = 32'hFFFFFFF1;
    // rom_array[37695] = 32'hFFFFFFF1;
    // rom_array[37696] = 32'hFFFFFFF1;
    // rom_array[37697] = 32'hFFFFFFF0;
    // rom_array[37698] = 32'hFFFFFFF0;
    // rom_array[37699] = 32'hFFFFFFF0;
    // rom_array[37700] = 32'hFFFFFFF0;
    // rom_array[37701] = 32'hFFFFFFF1;
    // rom_array[37702] = 32'hFFFFFFF1;
    // rom_array[37703] = 32'hFFFFFFF1;
    // rom_array[37704] = 32'hFFFFFFF1;
    // rom_array[37705] = 32'hFFFFFFF1;
    // rom_array[37706] = 32'hFFFFFFF1;
    // rom_array[37707] = 32'hFFFFFFF1;
    // rom_array[37708] = 32'hFFFFFFF1;
    // rom_array[37709] = 32'hFFFFFFF1;
    // rom_array[37710] = 32'hFFFFFFF1;
    // rom_array[37711] = 32'hFFFFFFF1;
    // rom_array[37712] = 32'hFFFFFFF1;
    // rom_array[37713] = 32'hFFFFFFF1;
    // rom_array[37714] = 32'hFFFFFFF1;
    // rom_array[37715] = 32'hFFFFFFF1;
    // rom_array[37716] = 32'hFFFFFFF1;
    // rom_array[37717] = 32'hFFFFFFF1;
    // rom_array[37718] = 32'hFFFFFFF1;
    // rom_array[37719] = 32'hFFFFFFF1;
    // rom_array[37720] = 32'hFFFFFFF1;
    // rom_array[37721] = 32'hFFFFFFF0;
    // rom_array[37722] = 32'hFFFFFFF0;
    // rom_array[37723] = 32'hFFFFFFF0;
    // rom_array[37724] = 32'hFFFFFFF0;
    // rom_array[37725] = 32'hFFFFFFF1;
    // rom_array[37726] = 32'hFFFFFFF1;
    // rom_array[37727] = 32'hFFFFFFF1;
    // rom_array[37728] = 32'hFFFFFFF1;
    // rom_array[37729] = 32'hFFFFFFF0;
    // rom_array[37730] = 32'hFFFFFFF0;
    // rom_array[37731] = 32'hFFFFFFF0;
    // rom_array[37732] = 32'hFFFFFFF0;
    // rom_array[37733] = 32'hFFFFFFF1;
    // rom_array[37734] = 32'hFFFFFFF1;
    // rom_array[37735] = 32'hFFFFFFF1;
    // rom_array[37736] = 32'hFFFFFFF1;
    // rom_array[37737] = 32'hFFFFFFF0;
    // rom_array[37738] = 32'hFFFFFFF0;
    // rom_array[37739] = 32'hFFFFFFF0;
    // rom_array[37740] = 32'hFFFFFFF0;
    // rom_array[37741] = 32'hFFFFFFF1;
    // rom_array[37742] = 32'hFFFFFFF1;
    // rom_array[37743] = 32'hFFFFFFF1;
    // rom_array[37744] = 32'hFFFFFFF1;
    // rom_array[37745] = 32'hFFFFFFF0;
    // rom_array[37746] = 32'hFFFFFFF0;
    // rom_array[37747] = 32'hFFFFFFF0;
    // rom_array[37748] = 32'hFFFFFFF0;
    // rom_array[37749] = 32'hFFFFFFF1;
    // rom_array[37750] = 32'hFFFFFFF1;
    // rom_array[37751] = 32'hFFFFFFF1;
    // rom_array[37752] = 32'hFFFFFFF1;
    // rom_array[37753] = 32'hFFFFFFF1;
    // rom_array[37754] = 32'hFFFFFFF1;
    // rom_array[37755] = 32'hFFFFFFF1;
    // rom_array[37756] = 32'hFFFFFFF1;
    // rom_array[37757] = 32'hFFFFFFF1;
    // rom_array[37758] = 32'hFFFFFFF1;
    // rom_array[37759] = 32'hFFFFFFF1;
    // rom_array[37760] = 32'hFFFFFFF1;
    // rom_array[37761] = 32'hFFFFFFF1;
    // rom_array[37762] = 32'hFFFFFFF1;
    // rom_array[37763] = 32'hFFFFFFF1;
    // rom_array[37764] = 32'hFFFFFFF1;
    // rom_array[37765] = 32'hFFFFFFF1;
    // rom_array[37766] = 32'hFFFFFFF1;
    // rom_array[37767] = 32'hFFFFFFF1;
    // rom_array[37768] = 32'hFFFFFFF1;
    // rom_array[37769] = 32'hFFFFFFF1;
    // rom_array[37770] = 32'hFFFFFFF1;
    // rom_array[37771] = 32'hFFFFFFF1;
    // rom_array[37772] = 32'hFFFFFFF1;
    // rom_array[37773] = 32'hFFFFFFF1;
    // rom_array[37774] = 32'hFFFFFFF1;
    // rom_array[37775] = 32'hFFFFFFF1;
    // rom_array[37776] = 32'hFFFFFFF1;
    // rom_array[37777] = 32'hFFFFFFF1;
    // rom_array[37778] = 32'hFFFFFFF1;
    // rom_array[37779] = 32'hFFFFFFF1;
    // rom_array[37780] = 32'hFFFFFFF1;
    // rom_array[37781] = 32'hFFFFFFF1;
    // rom_array[37782] = 32'hFFFFFFF1;
    // rom_array[37783] = 32'hFFFFFFF1;
    // rom_array[37784] = 32'hFFFFFFF1;
    // rom_array[37785] = 32'hFFFFFFF1;
    // rom_array[37786] = 32'hFFFFFFF1;
    // rom_array[37787] = 32'hFFFFFFF1;
    // rom_array[37788] = 32'hFFFFFFF1;
    // rom_array[37789] = 32'hFFFFFFF0;
    // rom_array[37790] = 32'hFFFFFFF0;
    // rom_array[37791] = 32'hFFFFFFF1;
    // rom_array[37792] = 32'hFFFFFFF1;
    // rom_array[37793] = 32'hFFFFFFF1;
    // rom_array[37794] = 32'hFFFFFFF1;
    // rom_array[37795] = 32'hFFFFFFF1;
    // rom_array[37796] = 32'hFFFFFFF1;
    // rom_array[37797] = 32'hFFFFFFF0;
    // rom_array[37798] = 32'hFFFFFFF0;
    // rom_array[37799] = 32'hFFFFFFF1;
    // rom_array[37800] = 32'hFFFFFFF1;
    // rom_array[37801] = 32'hFFFFFFF1;
    // rom_array[37802] = 32'hFFFFFFF1;
    // rom_array[37803] = 32'hFFFFFFF1;
    // rom_array[37804] = 32'hFFFFFFF1;
    // rom_array[37805] = 32'hFFFFFFF0;
    // rom_array[37806] = 32'hFFFFFFF0;
    // rom_array[37807] = 32'hFFFFFFF0;
    // rom_array[37808] = 32'hFFFFFFF0;
    // rom_array[37809] = 32'hFFFFFFF1;
    // rom_array[37810] = 32'hFFFFFFF1;
    // rom_array[37811] = 32'hFFFFFFF1;
    // rom_array[37812] = 32'hFFFFFFF1;
    // rom_array[37813] = 32'hFFFFFFF0;
    // rom_array[37814] = 32'hFFFFFFF0;
    // rom_array[37815] = 32'hFFFFFFF0;
    // rom_array[37816] = 32'hFFFFFFF0;
    // rom_array[37817] = 32'hFFFFFFF0;
    // rom_array[37818] = 32'hFFFFFFF0;
    // rom_array[37819] = 32'hFFFFFFF1;
    // rom_array[37820] = 32'hFFFFFFF1;
    // rom_array[37821] = 32'hFFFFFFF0;
    // rom_array[37822] = 32'hFFFFFFF0;
    // rom_array[37823] = 32'hFFFFFFF1;
    // rom_array[37824] = 32'hFFFFFFF1;
    // rom_array[37825] = 32'hFFFFFFF0;
    // rom_array[37826] = 32'hFFFFFFF0;
    // rom_array[37827] = 32'hFFFFFFF1;
    // rom_array[37828] = 32'hFFFFFFF1;
    // rom_array[37829] = 32'hFFFFFFF0;
    // rom_array[37830] = 32'hFFFFFFF0;
    // rom_array[37831] = 32'hFFFFFFF1;
    // rom_array[37832] = 32'hFFFFFFF1;
    // rom_array[37833] = 32'hFFFFFFF1;
    // rom_array[37834] = 32'hFFFFFFF1;
    // rom_array[37835] = 32'hFFFFFFF1;
    // rom_array[37836] = 32'hFFFFFFF1;
    // rom_array[37837] = 32'hFFFFFFF0;
    // rom_array[37838] = 32'hFFFFFFF0;
    // rom_array[37839] = 32'hFFFFFFF0;
    // rom_array[37840] = 32'hFFFFFFF0;
    // rom_array[37841] = 32'hFFFFFFF1;
    // rom_array[37842] = 32'hFFFFFFF1;
    // rom_array[37843] = 32'hFFFFFFF1;
    // rom_array[37844] = 32'hFFFFFFF1;
    // rom_array[37845] = 32'hFFFFFFF0;
    // rom_array[37846] = 32'hFFFFFFF0;
    // rom_array[37847] = 32'hFFFFFFF0;
    // rom_array[37848] = 32'hFFFFFFF0;
    // rom_array[37849] = 32'hFFFFFFF1;
    // rom_array[37850] = 32'hFFFFFFF1;
    // rom_array[37851] = 32'hFFFFFFF1;
    // rom_array[37852] = 32'hFFFFFFF1;
    // rom_array[37853] = 32'hFFFFFFF0;
    // rom_array[37854] = 32'hFFFFFFF0;
    // rom_array[37855] = 32'hFFFFFFF0;
    // rom_array[37856] = 32'hFFFFFFF0;
    // rom_array[37857] = 32'hFFFFFFF1;
    // rom_array[37858] = 32'hFFFFFFF1;
    // rom_array[37859] = 32'hFFFFFFF1;
    // rom_array[37860] = 32'hFFFFFFF1;
    // rom_array[37861] = 32'hFFFFFFF0;
    // rom_array[37862] = 32'hFFFFFFF0;
    // rom_array[37863] = 32'hFFFFFFF0;
    // rom_array[37864] = 32'hFFFFFFF0;
    // rom_array[37865] = 32'hFFFFFFF0;
    // rom_array[37866] = 32'hFFFFFFF0;
    // rom_array[37867] = 32'hFFFFFFF1;
    // rom_array[37868] = 32'hFFFFFFF1;
    // rom_array[37869] = 32'hFFFFFFF0;
    // rom_array[37870] = 32'hFFFFFFF0;
    // rom_array[37871] = 32'hFFFFFFF1;
    // rom_array[37872] = 32'hFFFFFFF1;
    // rom_array[37873] = 32'hFFFFFFF0;
    // rom_array[37874] = 32'hFFFFFFF0;
    // rom_array[37875] = 32'hFFFFFFF1;
    // rom_array[37876] = 32'hFFFFFFF1;
    // rom_array[37877] = 32'hFFFFFFF0;
    // rom_array[37878] = 32'hFFFFFFF0;
    // rom_array[37879] = 32'hFFFFFFF1;
    // rom_array[37880] = 32'hFFFFFFF1;
    // rom_array[37881] = 32'hFFFFFFF0;
    // rom_array[37882] = 32'hFFFFFFF0;
    // rom_array[37883] = 32'hFFFFFFF1;
    // rom_array[37884] = 32'hFFFFFFF1;
    // rom_array[37885] = 32'hFFFFFFF0;
    // rom_array[37886] = 32'hFFFFFFF0;
    // rom_array[37887] = 32'hFFFFFFF0;
    // rom_array[37888] = 32'hFFFFFFF0;
    // rom_array[37889] = 32'hFFFFFFF0;
    // rom_array[37890] = 32'hFFFFFFF0;
    // rom_array[37891] = 32'hFFFFFFF1;
    // rom_array[37892] = 32'hFFFFFFF1;
    // rom_array[37893] = 32'hFFFFFFF0;
    // rom_array[37894] = 32'hFFFFFFF0;
    // rom_array[37895] = 32'hFFFFFFF0;
    // rom_array[37896] = 32'hFFFFFFF0;
    // rom_array[37897] = 32'hFFFFFFF1;
    // rom_array[37898] = 32'hFFFFFFF1;
    // rom_array[37899] = 32'hFFFFFFF1;
    // rom_array[37900] = 32'hFFFFFFF1;
    // rom_array[37901] = 32'hFFFFFFF0;
    // rom_array[37902] = 32'hFFFFFFF0;
    // rom_array[37903] = 32'hFFFFFFF0;
    // rom_array[37904] = 32'hFFFFFFF0;
    // rom_array[37905] = 32'hFFFFFFF1;
    // rom_array[37906] = 32'hFFFFFFF1;
    // rom_array[37907] = 32'hFFFFFFF1;
    // rom_array[37908] = 32'hFFFFFFF1;
    // rom_array[37909] = 32'hFFFFFFF0;
    // rom_array[37910] = 32'hFFFFFFF0;
    // rom_array[37911] = 32'hFFFFFFF0;
    // rom_array[37912] = 32'hFFFFFFF0;
    // rom_array[37913] = 32'hFFFFFFF1;
    // rom_array[37914] = 32'hFFFFFFF1;
    // rom_array[37915] = 32'hFFFFFFF1;
    // rom_array[37916] = 32'hFFFFFFF1;
    // rom_array[37917] = 32'hFFFFFFF0;
    // rom_array[37918] = 32'hFFFFFFF0;
    // rom_array[37919] = 32'hFFFFFFF0;
    // rom_array[37920] = 32'hFFFFFFF0;
    // rom_array[37921] = 32'hFFFFFFF1;
    // rom_array[37922] = 32'hFFFFFFF1;
    // rom_array[37923] = 32'hFFFFFFF1;
    // rom_array[37924] = 32'hFFFFFFF1;
    // rom_array[37925] = 32'hFFFFFFF0;
    // rom_array[37926] = 32'hFFFFFFF0;
    // rom_array[37927] = 32'hFFFFFFF0;
    // rom_array[37928] = 32'hFFFFFFF0;
    // rom_array[37929] = 32'hFFFFFFF1;
    // rom_array[37930] = 32'hFFFFFFF1;
    // rom_array[37931] = 32'hFFFFFFF1;
    // rom_array[37932] = 32'hFFFFFFF1;
    // rom_array[37933] = 32'hFFFFFFF0;
    // rom_array[37934] = 32'hFFFFFFF0;
    // rom_array[37935] = 32'hFFFFFFF0;
    // rom_array[37936] = 32'hFFFFFFF0;
    // rom_array[37937] = 32'hFFFFFFF1;
    // rom_array[37938] = 32'hFFFFFFF1;
    // rom_array[37939] = 32'hFFFFFFF1;
    // rom_array[37940] = 32'hFFFFFFF1;
    // rom_array[37941] = 32'hFFFFFFF0;
    // rom_array[37942] = 32'hFFFFFFF0;
    // rom_array[37943] = 32'hFFFFFFF0;
    // rom_array[37944] = 32'hFFFFFFF0;
    // rom_array[37945] = 32'hFFFFFFF1;
    // rom_array[37946] = 32'hFFFFFFF1;
    // rom_array[37947] = 32'hFFFFFFF1;
    // rom_array[37948] = 32'hFFFFFFF1;
    // rom_array[37949] = 32'hFFFFFFF1;
    // rom_array[37950] = 32'hFFFFFFF1;
    // rom_array[37951] = 32'hFFFFFFF1;
    // rom_array[37952] = 32'hFFFFFFF1;
    // rom_array[37953] = 32'hFFFFFFF1;
    // rom_array[37954] = 32'hFFFFFFF1;
    // rom_array[37955] = 32'hFFFFFFF1;
    // rom_array[37956] = 32'hFFFFFFF1;
    // rom_array[37957] = 32'hFFFFFFF1;
    // rom_array[37958] = 32'hFFFFFFF1;
    // rom_array[37959] = 32'hFFFFFFF1;
    // rom_array[37960] = 32'hFFFFFFF1;
    // rom_array[37961] = 32'hFFFFFFF1;
    // rom_array[37962] = 32'hFFFFFFF1;
    // rom_array[37963] = 32'hFFFFFFF1;
    // rom_array[37964] = 32'hFFFFFFF1;
    // rom_array[37965] = 32'hFFFFFFF0;
    // rom_array[37966] = 32'hFFFFFFF0;
    // rom_array[37967] = 32'hFFFFFFF0;
    // rom_array[37968] = 32'hFFFFFFF0;
    // rom_array[37969] = 32'hFFFFFFF1;
    // rom_array[37970] = 32'hFFFFFFF1;
    // rom_array[37971] = 32'hFFFFFFF1;
    // rom_array[37972] = 32'hFFFFFFF1;
    // rom_array[37973] = 32'hFFFFFFF0;
    // rom_array[37974] = 32'hFFFFFFF0;
    // rom_array[37975] = 32'hFFFFFFF0;
    // rom_array[37976] = 32'hFFFFFFF0;
    // rom_array[37977] = 32'hFFFFFFF1;
    // rom_array[37978] = 32'hFFFFFFF1;
    // rom_array[37979] = 32'hFFFFFFF1;
    // rom_array[37980] = 32'hFFFFFFF1;
    // rom_array[37981] = 32'hFFFFFFF1;
    // rom_array[37982] = 32'hFFFFFFF1;
    // rom_array[37983] = 32'hFFFFFFF1;
    // rom_array[37984] = 32'hFFFFFFF1;
    // rom_array[37985] = 32'hFFFFFFF1;
    // rom_array[37986] = 32'hFFFFFFF1;
    // rom_array[37987] = 32'hFFFFFFF1;
    // rom_array[37988] = 32'hFFFFFFF1;
    // rom_array[37989] = 32'hFFFFFFF1;
    // rom_array[37990] = 32'hFFFFFFF1;
    // rom_array[37991] = 32'hFFFFFFF1;
    // rom_array[37992] = 32'hFFFFFFF1;
    // rom_array[37993] = 32'hFFFFFFF1;
    // rom_array[37994] = 32'hFFFFFFF1;
    // rom_array[37995] = 32'hFFFFFFF1;
    // rom_array[37996] = 32'hFFFFFFF1;
    // rom_array[37997] = 32'hFFFFFFF0;
    // rom_array[37998] = 32'hFFFFFFF0;
    // rom_array[37999] = 32'hFFFFFFF0;
    // rom_array[38000] = 32'hFFFFFFF0;
    // rom_array[38001] = 32'hFFFFFFF1;
    // rom_array[38002] = 32'hFFFFFFF1;
    // rom_array[38003] = 32'hFFFFFFF1;
    // rom_array[38004] = 32'hFFFFFFF1;
    // rom_array[38005] = 32'hFFFFFFF0;
    // rom_array[38006] = 32'hFFFFFFF0;
    // rom_array[38007] = 32'hFFFFFFF0;
    // rom_array[38008] = 32'hFFFFFFF0;
    // rom_array[38009] = 32'hFFFFFFF1;
    // rom_array[38010] = 32'hFFFFFFF1;
    // rom_array[38011] = 32'hFFFFFFF1;
    // rom_array[38012] = 32'hFFFFFFF1;
    // rom_array[38013] = 32'hFFFFFFF0;
    // rom_array[38014] = 32'hFFFFFFF0;
    // rom_array[38015] = 32'hFFFFFFF0;
    // rom_array[38016] = 32'hFFFFFFF0;
    // rom_array[38017] = 32'hFFFFFFF1;
    // rom_array[38018] = 32'hFFFFFFF1;
    // rom_array[38019] = 32'hFFFFFFF1;
    // rom_array[38020] = 32'hFFFFFFF1;
    // rom_array[38021] = 32'hFFFFFFF0;
    // rom_array[38022] = 32'hFFFFFFF0;
    // rom_array[38023] = 32'hFFFFFFF0;
    // rom_array[38024] = 32'hFFFFFFF0;
    // rom_array[38025] = 32'hFFFFFFF1;
    // rom_array[38026] = 32'hFFFFFFF1;
    // rom_array[38027] = 32'hFFFFFFF1;
    // rom_array[38028] = 32'hFFFFFFF1;
    // rom_array[38029] = 32'hFFFFFFF1;
    // rom_array[38030] = 32'hFFFFFFF1;
    // rom_array[38031] = 32'hFFFFFFF1;
    // rom_array[38032] = 32'hFFFFFFF1;
    // rom_array[38033] = 32'hFFFFFFF1;
    // rom_array[38034] = 32'hFFFFFFF1;
    // rom_array[38035] = 32'hFFFFFFF1;
    // rom_array[38036] = 32'hFFFFFFF1;
    // rom_array[38037] = 32'hFFFFFFF1;
    // rom_array[38038] = 32'hFFFFFFF1;
    // rom_array[38039] = 32'hFFFFFFF1;
    // rom_array[38040] = 32'hFFFFFFF1;
    // rom_array[38041] = 32'hFFFFFFF1;
    // rom_array[38042] = 32'hFFFFFFF1;
    // rom_array[38043] = 32'hFFFFFFF1;
    // rom_array[38044] = 32'hFFFFFFF1;
    // rom_array[38045] = 32'hFFFFFFF0;
    // rom_array[38046] = 32'hFFFFFFF0;
    // rom_array[38047] = 32'hFFFFFFF0;
    // rom_array[38048] = 32'hFFFFFFF0;
    // rom_array[38049] = 32'hFFFFFFF1;
    // rom_array[38050] = 32'hFFFFFFF1;
    // rom_array[38051] = 32'hFFFFFFF1;
    // rom_array[38052] = 32'hFFFFFFF1;
    // rom_array[38053] = 32'hFFFFFFF0;
    // rom_array[38054] = 32'hFFFFFFF0;
    // rom_array[38055] = 32'hFFFFFFF0;
    // rom_array[38056] = 32'hFFFFFFF0;
    // rom_array[38057] = 32'hFFFFFFF0;
    // rom_array[38058] = 32'hFFFFFFF0;
    // rom_array[38059] = 32'hFFFFFFF1;
    // rom_array[38060] = 32'hFFFFFFF1;
    // rom_array[38061] = 32'hFFFFFFF0;
    // rom_array[38062] = 32'hFFFFFFF0;
    // rom_array[38063] = 32'hFFFFFFF1;
    // rom_array[38064] = 32'hFFFFFFF1;
    // rom_array[38065] = 32'hFFFFFFF0;
    // rom_array[38066] = 32'hFFFFFFF0;
    // rom_array[38067] = 32'hFFFFFFF1;
    // rom_array[38068] = 32'hFFFFFFF1;
    // rom_array[38069] = 32'hFFFFFFF0;
    // rom_array[38070] = 32'hFFFFFFF0;
    // rom_array[38071] = 32'hFFFFFFF1;
    // rom_array[38072] = 32'hFFFFFFF1;
    // rom_array[38073] = 32'hFFFFFFF1;
    // rom_array[38074] = 32'hFFFFFFF1;
    // rom_array[38075] = 32'hFFFFFFF1;
    // rom_array[38076] = 32'hFFFFFFF1;
    // rom_array[38077] = 32'hFFFFFFF1;
    // rom_array[38078] = 32'hFFFFFFF1;
    // rom_array[38079] = 32'hFFFFFFF1;
    // rom_array[38080] = 32'hFFFFFFF1;
    // rom_array[38081] = 32'hFFFFFFF1;
    // rom_array[38082] = 32'hFFFFFFF1;
    // rom_array[38083] = 32'hFFFFFFF1;
    // rom_array[38084] = 32'hFFFFFFF1;
    // rom_array[38085] = 32'hFFFFFFF1;
    // rom_array[38086] = 32'hFFFFFFF1;
    // rom_array[38087] = 32'hFFFFFFF1;
    // rom_array[38088] = 32'hFFFFFFF1;
    // rom_array[38089] = 32'hFFFFFFF0;
    // rom_array[38090] = 32'hFFFFFFF0;
    // rom_array[38091] = 32'hFFFFFFF1;
    // rom_array[38092] = 32'hFFFFFFF1;
    // rom_array[38093] = 32'hFFFFFFF0;
    // rom_array[38094] = 32'hFFFFFFF0;
    // rom_array[38095] = 32'hFFFFFFF1;
    // rom_array[38096] = 32'hFFFFFFF1;
    // rom_array[38097] = 32'hFFFFFFF0;
    // rom_array[38098] = 32'hFFFFFFF0;
    // rom_array[38099] = 32'hFFFFFFF1;
    // rom_array[38100] = 32'hFFFFFFF1;
    // rom_array[38101] = 32'hFFFFFFF0;
    // rom_array[38102] = 32'hFFFFFFF0;
    // rom_array[38103] = 32'hFFFFFFF1;
    // rom_array[38104] = 32'hFFFFFFF1;
    // rom_array[38105] = 32'hFFFFFFF1;
    // rom_array[38106] = 32'hFFFFFFF1;
    // rom_array[38107] = 32'hFFFFFFF1;
    // rom_array[38108] = 32'hFFFFFFF1;
    // rom_array[38109] = 32'hFFFFFFF1;
    // rom_array[38110] = 32'hFFFFFFF1;
    // rom_array[38111] = 32'hFFFFFFF1;
    // rom_array[38112] = 32'hFFFFFFF1;
    // rom_array[38113] = 32'hFFFFFFF1;
    // rom_array[38114] = 32'hFFFFFFF1;
    // rom_array[38115] = 32'hFFFFFFF1;
    // rom_array[38116] = 32'hFFFFFFF1;
    // rom_array[38117] = 32'hFFFFFFF1;
    // rom_array[38118] = 32'hFFFFFFF1;
    // rom_array[38119] = 32'hFFFFFFF1;
    // rom_array[38120] = 32'hFFFFFFF1;
    // rom_array[38121] = 32'hFFFFFFF1;
    // rom_array[38122] = 32'hFFFFFFF1;
    // rom_array[38123] = 32'hFFFFFFF1;
    // rom_array[38124] = 32'hFFFFFFF1;
    // rom_array[38125] = 32'hFFFFFFF1;
    // rom_array[38126] = 32'hFFFFFFF1;
    // rom_array[38127] = 32'hFFFFFFF1;
    // rom_array[38128] = 32'hFFFFFFF1;
    // rom_array[38129] = 32'hFFFFFFF1;
    // rom_array[38130] = 32'hFFFFFFF1;
    // rom_array[38131] = 32'hFFFFFFF1;
    // rom_array[38132] = 32'hFFFFFFF1;
    // rom_array[38133] = 32'hFFFFFFF1;
    // rom_array[38134] = 32'hFFFFFFF1;
    // rom_array[38135] = 32'hFFFFFFF1;
    // rom_array[38136] = 32'hFFFFFFF1;
    // rom_array[38137] = 32'hFFFFFFF1;
    // rom_array[38138] = 32'hFFFFFFF1;
    // rom_array[38139] = 32'hFFFFFFF1;
    // rom_array[38140] = 32'hFFFFFFF1;
    // rom_array[38141] = 32'hFFFFFFF1;
    // rom_array[38142] = 32'hFFFFFFF1;
    // rom_array[38143] = 32'hFFFFFFF1;
    // rom_array[38144] = 32'hFFFFFFF1;
    // rom_array[38145] = 32'hFFFFFFF1;
    // rom_array[38146] = 32'hFFFFFFF1;
    // rom_array[38147] = 32'hFFFFFFF1;
    // rom_array[38148] = 32'hFFFFFFF1;
    // rom_array[38149] = 32'hFFFFFFF1;
    // rom_array[38150] = 32'hFFFFFFF1;
    // rom_array[38151] = 32'hFFFFFFF1;
    // rom_array[38152] = 32'hFFFFFFF1;
    // rom_array[38153] = 32'hFFFFFFF0;
    // rom_array[38154] = 32'hFFFFFFF0;
    // rom_array[38155] = 32'hFFFFFFF1;
    // rom_array[38156] = 32'hFFFFFFF1;
    // rom_array[38157] = 32'hFFFFFFF0;
    // rom_array[38158] = 32'hFFFFFFF0;
    // rom_array[38159] = 32'hFFFFFFF1;
    // rom_array[38160] = 32'hFFFFFFF1;
    // rom_array[38161] = 32'hFFFFFFF0;
    // rom_array[38162] = 32'hFFFFFFF0;
    // rom_array[38163] = 32'hFFFFFFF1;
    // rom_array[38164] = 32'hFFFFFFF1;
    // rom_array[38165] = 32'hFFFFFFF0;
    // rom_array[38166] = 32'hFFFFFFF0;
    // rom_array[38167] = 32'hFFFFFFF1;
    // rom_array[38168] = 32'hFFFFFFF1;
    // rom_array[38169] = 32'hFFFFFFF0;
    // rom_array[38170] = 32'hFFFFFFF0;
    // rom_array[38171] = 32'hFFFFFFF1;
    // rom_array[38172] = 32'hFFFFFFF1;
    // rom_array[38173] = 32'hFFFFFFF0;
    // rom_array[38174] = 32'hFFFFFFF0;
    // rom_array[38175] = 32'hFFFFFFF1;
    // rom_array[38176] = 32'hFFFFFFF1;
    // rom_array[38177] = 32'hFFFFFFF0;
    // rom_array[38178] = 32'hFFFFFFF0;
    // rom_array[38179] = 32'hFFFFFFF1;
    // rom_array[38180] = 32'hFFFFFFF1;
    // rom_array[38181] = 32'hFFFFFFF0;
    // rom_array[38182] = 32'hFFFFFFF0;
    // rom_array[38183] = 32'hFFFFFFF1;
    // rom_array[38184] = 32'hFFFFFFF1;
    // rom_array[38185] = 32'hFFFFFFF1;
    // rom_array[38186] = 32'hFFFFFFF1;
    // rom_array[38187] = 32'hFFFFFFF1;
    // rom_array[38188] = 32'hFFFFFFF1;
    // rom_array[38189] = 32'hFFFFFFF0;
    // rom_array[38190] = 32'hFFFFFFF0;
    // rom_array[38191] = 32'hFFFFFFF0;
    // rom_array[38192] = 32'hFFFFFFF0;
    // rom_array[38193] = 32'hFFFFFFF1;
    // rom_array[38194] = 32'hFFFFFFF1;
    // rom_array[38195] = 32'hFFFFFFF1;
    // rom_array[38196] = 32'hFFFFFFF1;
    // rom_array[38197] = 32'hFFFFFFF0;
    // rom_array[38198] = 32'hFFFFFFF0;
    // rom_array[38199] = 32'hFFFFFFF0;
    // rom_array[38200] = 32'hFFFFFFF0;
    // rom_array[38201] = 32'hFFFFFFF1;
    // rom_array[38202] = 32'hFFFFFFF1;
    // rom_array[38203] = 32'hFFFFFFF1;
    // rom_array[38204] = 32'hFFFFFFF1;
    // rom_array[38205] = 32'hFFFFFFF1;
    // rom_array[38206] = 32'hFFFFFFF1;
    // rom_array[38207] = 32'hFFFFFFF1;
    // rom_array[38208] = 32'hFFFFFFF1;
    // rom_array[38209] = 32'hFFFFFFF1;
    // rom_array[38210] = 32'hFFFFFFF1;
    // rom_array[38211] = 32'hFFFFFFF1;
    // rom_array[38212] = 32'hFFFFFFF1;
    // rom_array[38213] = 32'hFFFFFFF1;
    // rom_array[38214] = 32'hFFFFFFF1;
    // rom_array[38215] = 32'hFFFFFFF1;
    // rom_array[38216] = 32'hFFFFFFF1;
    // rom_array[38217] = 32'hFFFFFFF1;
    // rom_array[38218] = 32'hFFFFFFF1;
    // rom_array[38219] = 32'hFFFFFFF1;
    // rom_array[38220] = 32'hFFFFFFF1;
    // rom_array[38221] = 32'hFFFFFFF1;
    // rom_array[38222] = 32'hFFFFFFF1;
    // rom_array[38223] = 32'hFFFFFFF0;
    // rom_array[38224] = 32'hFFFFFFF0;
    // rom_array[38225] = 32'hFFFFFFF1;
    // rom_array[38226] = 32'hFFFFFFF1;
    // rom_array[38227] = 32'hFFFFFFF1;
    // rom_array[38228] = 32'hFFFFFFF1;
    // rom_array[38229] = 32'hFFFFFFF1;
    // rom_array[38230] = 32'hFFFFFFF1;
    // rom_array[38231] = 32'hFFFFFFF0;
    // rom_array[38232] = 32'hFFFFFFF0;
    // rom_array[38233] = 32'hFFFFFFF0;
    // rom_array[38234] = 32'hFFFFFFF0;
    // rom_array[38235] = 32'hFFFFFFF1;
    // rom_array[38236] = 32'hFFFFFFF1;
    // rom_array[38237] = 32'hFFFFFFF0;
    // rom_array[38238] = 32'hFFFFFFF0;
    // rom_array[38239] = 32'hFFFFFFF0;
    // rom_array[38240] = 32'hFFFFFFF0;
    // rom_array[38241] = 32'hFFFFFFF0;
    // rom_array[38242] = 32'hFFFFFFF0;
    // rom_array[38243] = 32'hFFFFFFF1;
    // rom_array[38244] = 32'hFFFFFFF1;
    // rom_array[38245] = 32'hFFFFFFF0;
    // rom_array[38246] = 32'hFFFFFFF0;
    // rom_array[38247] = 32'hFFFFFFF0;
    // rom_array[38248] = 32'hFFFFFFF0;
    // rom_array[38249] = 32'hFFFFFFF1;
    // rom_array[38250] = 32'hFFFFFFF1;
    // rom_array[38251] = 32'hFFFFFFF1;
    // rom_array[38252] = 32'hFFFFFFF1;
    // rom_array[38253] = 32'hFFFFFFF0;
    // rom_array[38254] = 32'hFFFFFFF0;
    // rom_array[38255] = 32'hFFFFFFF0;
    // rom_array[38256] = 32'hFFFFFFF0;
    // rom_array[38257] = 32'hFFFFFFF1;
    // rom_array[38258] = 32'hFFFFFFF1;
    // rom_array[38259] = 32'hFFFFFFF1;
    // rom_array[38260] = 32'hFFFFFFF1;
    // rom_array[38261] = 32'hFFFFFFF0;
    // rom_array[38262] = 32'hFFFFFFF0;
    // rom_array[38263] = 32'hFFFFFFF0;
    // rom_array[38264] = 32'hFFFFFFF0;
    // rom_array[38265] = 32'hFFFFFFF1;
    // rom_array[38266] = 32'hFFFFFFF1;
    // rom_array[38267] = 32'hFFFFFFF1;
    // rom_array[38268] = 32'hFFFFFFF1;
    // rom_array[38269] = 32'hFFFFFFF0;
    // rom_array[38270] = 32'hFFFFFFF0;
    // rom_array[38271] = 32'hFFFFFFF0;
    // rom_array[38272] = 32'hFFFFFFF0;
    // rom_array[38273] = 32'hFFFFFFF1;
    // rom_array[38274] = 32'hFFFFFFF1;
    // rom_array[38275] = 32'hFFFFFFF1;
    // rom_array[38276] = 32'hFFFFFFF1;
    // rom_array[38277] = 32'hFFFFFFF0;
    // rom_array[38278] = 32'hFFFFFFF0;
    // rom_array[38279] = 32'hFFFFFFF0;
    // rom_array[38280] = 32'hFFFFFFF0;
    // rom_array[38281] = 32'hFFFFFFF1;
    // rom_array[38282] = 32'hFFFFFFF1;
    // rom_array[38283] = 32'hFFFFFFF1;
    // rom_array[38284] = 32'hFFFFFFF1;
    // rom_array[38285] = 32'hFFFFFFF0;
    // rom_array[38286] = 32'hFFFFFFF0;
    // rom_array[38287] = 32'hFFFFFFF0;
    // rom_array[38288] = 32'hFFFFFFF0;
    // rom_array[38289] = 32'hFFFFFFF1;
    // rom_array[38290] = 32'hFFFFFFF1;
    // rom_array[38291] = 32'hFFFFFFF1;
    // rom_array[38292] = 32'hFFFFFFF1;
    // rom_array[38293] = 32'hFFFFFFF0;
    // rom_array[38294] = 32'hFFFFFFF0;
    // rom_array[38295] = 32'hFFFFFFF0;
    // rom_array[38296] = 32'hFFFFFFF0;
    // rom_array[38297] = 32'hFFFFFFF1;
    // rom_array[38298] = 32'hFFFFFFF1;
    // rom_array[38299] = 32'hFFFFFFF1;
    // rom_array[38300] = 32'hFFFFFFF1;
    // rom_array[38301] = 32'hFFFFFFF0;
    // rom_array[38302] = 32'hFFFFFFF0;
    // rom_array[38303] = 32'hFFFFFFF0;
    // rom_array[38304] = 32'hFFFFFFF0;
    // rom_array[38305] = 32'hFFFFFFF1;
    // rom_array[38306] = 32'hFFFFFFF1;
    // rom_array[38307] = 32'hFFFFFFF1;
    // rom_array[38308] = 32'hFFFFFFF1;
    // rom_array[38309] = 32'hFFFFFFF0;
    // rom_array[38310] = 32'hFFFFFFF0;
    // rom_array[38311] = 32'hFFFFFFF0;
    // rom_array[38312] = 32'hFFFFFFF0;
    // rom_array[38313] = 32'hFFFFFFF1;
    // rom_array[38314] = 32'hFFFFFFF1;
    // rom_array[38315] = 32'hFFFFFFF1;
    // rom_array[38316] = 32'hFFFFFFF1;
    // rom_array[38317] = 32'hFFFFFFF0;
    // rom_array[38318] = 32'hFFFFFFF0;
    // rom_array[38319] = 32'hFFFFFFF0;
    // rom_array[38320] = 32'hFFFFFFF0;
    // rom_array[38321] = 32'hFFFFFFF1;
    // rom_array[38322] = 32'hFFFFFFF1;
    // rom_array[38323] = 32'hFFFFFFF1;
    // rom_array[38324] = 32'hFFFFFFF1;
    // rom_array[38325] = 32'hFFFFFFF0;
    // rom_array[38326] = 32'hFFFFFFF0;
    // rom_array[38327] = 32'hFFFFFFF0;
    // rom_array[38328] = 32'hFFFFFFF0;
    // rom_array[38329] = 32'hFFFFFFF1;
    // rom_array[38330] = 32'hFFFFFFF1;
    // rom_array[38331] = 32'hFFFFFFF1;
    // rom_array[38332] = 32'hFFFFFFF1;
    // rom_array[38333] = 32'hFFFFFFF0;
    // rom_array[38334] = 32'hFFFFFFF0;
    // rom_array[38335] = 32'hFFFFFFF0;
    // rom_array[38336] = 32'hFFFFFFF0;
    // rom_array[38337] = 32'hFFFFFFF1;
    // rom_array[38338] = 32'hFFFFFFF1;
    // rom_array[38339] = 32'hFFFFFFF1;
    // rom_array[38340] = 32'hFFFFFFF1;
    // rom_array[38341] = 32'hFFFFFFF0;
    // rom_array[38342] = 32'hFFFFFFF0;
    // rom_array[38343] = 32'hFFFFFFF0;
    // rom_array[38344] = 32'hFFFFFFF0;
    // rom_array[38345] = 32'hFFFFFFF1;
    // rom_array[38346] = 32'hFFFFFFF1;
    // rom_array[38347] = 32'hFFFFFFF1;
    // rom_array[38348] = 32'hFFFFFFF1;
    // rom_array[38349] = 32'hFFFFFFF0;
    // rom_array[38350] = 32'hFFFFFFF0;
    // rom_array[38351] = 32'hFFFFFFF0;
    // rom_array[38352] = 32'hFFFFFFF0;
    // rom_array[38353] = 32'hFFFFFFF1;
    // rom_array[38354] = 32'hFFFFFFF1;
    // rom_array[38355] = 32'hFFFFFFF1;
    // rom_array[38356] = 32'hFFFFFFF1;
    // rom_array[38357] = 32'hFFFFFFF0;
    // rom_array[38358] = 32'hFFFFFFF0;
    // rom_array[38359] = 32'hFFFFFFF0;
    // rom_array[38360] = 32'hFFFFFFF0;
    // rom_array[38361] = 32'hFFFFFFF1;
    // rom_array[38362] = 32'hFFFFFFF1;
    // rom_array[38363] = 32'hFFFFFFF1;
    // rom_array[38364] = 32'hFFFFFFF1;
    // rom_array[38365] = 32'hFFFFFFF0;
    // rom_array[38366] = 32'hFFFFFFF0;
    // rom_array[38367] = 32'hFFFFFFF0;
    // rom_array[38368] = 32'hFFFFFFF0;
    // rom_array[38369] = 32'hFFFFFFF1;
    // rom_array[38370] = 32'hFFFFFFF1;
    // rom_array[38371] = 32'hFFFFFFF1;
    // rom_array[38372] = 32'hFFFFFFF1;
    // rom_array[38373] = 32'hFFFFFFF0;
    // rom_array[38374] = 32'hFFFFFFF0;
    // rom_array[38375] = 32'hFFFFFFF0;
    // rom_array[38376] = 32'hFFFFFFF0;
    // rom_array[38377] = 32'hFFFFFFF1;
    // rom_array[38378] = 32'hFFFFFFF1;
    // rom_array[38379] = 32'hFFFFFFF1;
    // rom_array[38380] = 32'hFFFFFFF1;
    // rom_array[38381] = 32'hFFFFFFF0;
    // rom_array[38382] = 32'hFFFFFFF0;
    // rom_array[38383] = 32'hFFFFFFF0;
    // rom_array[38384] = 32'hFFFFFFF0;
    // rom_array[38385] = 32'hFFFFFFF1;
    // rom_array[38386] = 32'hFFFFFFF1;
    // rom_array[38387] = 32'hFFFFFFF1;
    // rom_array[38388] = 32'hFFFFFFF1;
    // rom_array[38389] = 32'hFFFFFFF0;
    // rom_array[38390] = 32'hFFFFFFF0;
    // rom_array[38391] = 32'hFFFFFFF0;
    // rom_array[38392] = 32'hFFFFFFF0;
    // rom_array[38393] = 32'hFFFFFFF1;
    // rom_array[38394] = 32'hFFFFFFF1;
    // rom_array[38395] = 32'hFFFFFFF1;
    // rom_array[38396] = 32'hFFFFFFF1;
    // rom_array[38397] = 32'hFFFFFFF0;
    // rom_array[38398] = 32'hFFFFFFF0;
    // rom_array[38399] = 32'hFFFFFFF0;
    // rom_array[38400] = 32'hFFFFFFF0;
    // rom_array[38401] = 32'hFFFFFFF1;
    // rom_array[38402] = 32'hFFFFFFF1;
    // rom_array[38403] = 32'hFFFFFFF1;
    // rom_array[38404] = 32'hFFFFFFF1;
    // rom_array[38405] = 32'hFFFFFFF0;
    // rom_array[38406] = 32'hFFFFFFF0;
    // rom_array[38407] = 32'hFFFFFFF0;
    // rom_array[38408] = 32'hFFFFFFF0;
    // rom_array[38409] = 32'hFFFFFFF1;
    // rom_array[38410] = 32'hFFFFFFF1;
    // rom_array[38411] = 32'hFFFFFFF1;
    // rom_array[38412] = 32'hFFFFFFF1;
    // rom_array[38413] = 32'hFFFFFFF0;
    // rom_array[38414] = 32'hFFFFFFF0;
    // rom_array[38415] = 32'hFFFFFFF0;
    // rom_array[38416] = 32'hFFFFFFF0;
    // rom_array[38417] = 32'hFFFFFFF1;
    // rom_array[38418] = 32'hFFFFFFF1;
    // rom_array[38419] = 32'hFFFFFFF1;
    // rom_array[38420] = 32'hFFFFFFF1;
    // rom_array[38421] = 32'hFFFFFFF0;
    // rom_array[38422] = 32'hFFFFFFF0;
    // rom_array[38423] = 32'hFFFFFFF0;
    // rom_array[38424] = 32'hFFFFFFF0;
    // rom_array[38425] = 32'hFFFFFFF0;
    // rom_array[38426] = 32'hFFFFFFF0;
    // rom_array[38427] = 32'hFFFFFFF0;
    // rom_array[38428] = 32'hFFFFFFF0;
    // rom_array[38429] = 32'hFFFFFFF0;
    // rom_array[38430] = 32'hFFFFFFF0;
    // rom_array[38431] = 32'hFFFFFFF1;
    // rom_array[38432] = 32'hFFFFFFF1;
    // rom_array[38433] = 32'hFFFFFFF0;
    // rom_array[38434] = 32'hFFFFFFF0;
    // rom_array[38435] = 32'hFFFFFFF0;
    // rom_array[38436] = 32'hFFFFFFF0;
    // rom_array[38437] = 32'hFFFFFFF0;
    // rom_array[38438] = 32'hFFFFFFF0;
    // rom_array[38439] = 32'hFFFFFFF1;
    // rom_array[38440] = 32'hFFFFFFF1;
    // rom_array[38441] = 32'hFFFFFFF0;
    // rom_array[38442] = 32'hFFFFFFF0;
    // rom_array[38443] = 32'hFFFFFFF0;
    // rom_array[38444] = 32'hFFFFFFF0;
    // rom_array[38445] = 32'hFFFFFFF1;
    // rom_array[38446] = 32'hFFFFFFF1;
    // rom_array[38447] = 32'hFFFFFFF1;
    // rom_array[38448] = 32'hFFFFFFF1;
    // rom_array[38449] = 32'hFFFFFFF0;
    // rom_array[38450] = 32'hFFFFFFF0;
    // rom_array[38451] = 32'hFFFFFFF0;
    // rom_array[38452] = 32'hFFFFFFF0;
    // rom_array[38453] = 32'hFFFFFFF1;
    // rom_array[38454] = 32'hFFFFFFF1;
    // rom_array[38455] = 32'hFFFFFFF1;
    // rom_array[38456] = 32'hFFFFFFF1;
    // rom_array[38457] = 32'hFFFFFFF0;
    // rom_array[38458] = 32'hFFFFFFF0;
    // rom_array[38459] = 32'hFFFFFFF1;
    // rom_array[38460] = 32'hFFFFFFF1;
    // rom_array[38461] = 32'hFFFFFFF0;
    // rom_array[38462] = 32'hFFFFFFF0;
    // rom_array[38463] = 32'hFFFFFFF1;
    // rom_array[38464] = 32'hFFFFFFF1;
    // rom_array[38465] = 32'hFFFFFFF0;
    // rom_array[38466] = 32'hFFFFFFF0;
    // rom_array[38467] = 32'hFFFFFFF1;
    // rom_array[38468] = 32'hFFFFFFF1;
    // rom_array[38469] = 32'hFFFFFFF0;
    // rom_array[38470] = 32'hFFFFFFF0;
    // rom_array[38471] = 32'hFFFFFFF1;
    // rom_array[38472] = 32'hFFFFFFF1;
    // rom_array[38473] = 32'hFFFFFFF0;
    // rom_array[38474] = 32'hFFFFFFF0;
    // rom_array[38475] = 32'hFFFFFFF0;
    // rom_array[38476] = 32'hFFFFFFF0;
    // rom_array[38477] = 32'hFFFFFFF1;
    // rom_array[38478] = 32'hFFFFFFF1;
    // rom_array[38479] = 32'hFFFFFFF1;
    // rom_array[38480] = 32'hFFFFFFF1;
    // rom_array[38481] = 32'hFFFFFFF0;
    // rom_array[38482] = 32'hFFFFFFF0;
    // rom_array[38483] = 32'hFFFFFFF0;
    // rom_array[38484] = 32'hFFFFFFF0;
    // rom_array[38485] = 32'hFFFFFFF1;
    // rom_array[38486] = 32'hFFFFFFF1;
    // rom_array[38487] = 32'hFFFFFFF1;
    // rom_array[38488] = 32'hFFFFFFF1;
    // rom_array[38489] = 32'hFFFFFFF0;
    // rom_array[38490] = 32'hFFFFFFF0;
    // rom_array[38491] = 32'hFFFFFFF0;
    // rom_array[38492] = 32'hFFFFFFF0;
    // rom_array[38493] = 32'hFFFFFFF1;
    // rom_array[38494] = 32'hFFFFFFF1;
    // rom_array[38495] = 32'hFFFFFFF1;
    // rom_array[38496] = 32'hFFFFFFF1;
    // rom_array[38497] = 32'hFFFFFFF0;
    // rom_array[38498] = 32'hFFFFFFF0;
    // rom_array[38499] = 32'hFFFFFFF0;
    // rom_array[38500] = 32'hFFFFFFF0;
    // rom_array[38501] = 32'hFFFFFFF1;
    // rom_array[38502] = 32'hFFFFFFF1;
    // rom_array[38503] = 32'hFFFFFFF1;
    // rom_array[38504] = 32'hFFFFFFF1;
    // rom_array[38505] = 32'hFFFFFFF0;
    // rom_array[38506] = 32'hFFFFFFF0;
    // rom_array[38507] = 32'hFFFFFFF1;
    // rom_array[38508] = 32'hFFFFFFF1;
    // rom_array[38509] = 32'hFFFFFFF0;
    // rom_array[38510] = 32'hFFFFFFF0;
    // rom_array[38511] = 32'hFFFFFFF1;
    // rom_array[38512] = 32'hFFFFFFF1;
    // rom_array[38513] = 32'hFFFFFFF0;
    // rom_array[38514] = 32'hFFFFFFF0;
    // rom_array[38515] = 32'hFFFFFFF1;
    // rom_array[38516] = 32'hFFFFFFF1;
    // rom_array[38517] = 32'hFFFFFFF0;
    // rom_array[38518] = 32'hFFFFFFF0;
    // rom_array[38519] = 32'hFFFFFFF1;
    // rom_array[38520] = 32'hFFFFFFF1;
    // rom_array[38521] = 32'hFFFFFFF0;
    // rom_array[38522] = 32'hFFFFFFF0;
    // rom_array[38523] = 32'hFFFFFFF1;
    // rom_array[38524] = 32'hFFFFFFF1;
    // rom_array[38525] = 32'hFFFFFFF0;
    // rom_array[38526] = 32'hFFFFFFF0;
    // rom_array[38527] = 32'hFFFFFFF1;
    // rom_array[38528] = 32'hFFFFFFF1;
    // rom_array[38529] = 32'hFFFFFFF0;
    // rom_array[38530] = 32'hFFFFFFF0;
    // rom_array[38531] = 32'hFFFFFFF1;
    // rom_array[38532] = 32'hFFFFFFF1;
    // rom_array[38533] = 32'hFFFFFFF0;
    // rom_array[38534] = 32'hFFFFFFF0;
    // rom_array[38535] = 32'hFFFFFFF1;
    // rom_array[38536] = 32'hFFFFFFF1;
    // rom_array[38537] = 32'hFFFFFFF0;
    // rom_array[38538] = 32'hFFFFFFF0;
    // rom_array[38539] = 32'hFFFFFFF0;
    // rom_array[38540] = 32'hFFFFFFF0;
    // rom_array[38541] = 32'hFFFFFFF1;
    // rom_array[38542] = 32'hFFFFFFF1;
    // rom_array[38543] = 32'hFFFFFFF1;
    // rom_array[38544] = 32'hFFFFFFF1;
    // rom_array[38545] = 32'hFFFFFFF0;
    // rom_array[38546] = 32'hFFFFFFF0;
    // rom_array[38547] = 32'hFFFFFFF0;
    // rom_array[38548] = 32'hFFFFFFF0;
    // rom_array[38549] = 32'hFFFFFFF1;
    // rom_array[38550] = 32'hFFFFFFF1;
    // rom_array[38551] = 32'hFFFFFFF1;
    // rom_array[38552] = 32'hFFFFFFF1;
    // rom_array[38553] = 32'hFFFFFFF0;
    // rom_array[38554] = 32'hFFFFFFF0;
    // rom_array[38555] = 32'hFFFFFFF0;
    // rom_array[38556] = 32'hFFFFFFF0;
    // rom_array[38557] = 32'hFFFFFFF1;
    // rom_array[38558] = 32'hFFFFFFF1;
    // rom_array[38559] = 32'hFFFFFFF1;
    // rom_array[38560] = 32'hFFFFFFF1;
    // rom_array[38561] = 32'hFFFFFFF0;
    // rom_array[38562] = 32'hFFFFFFF0;
    // rom_array[38563] = 32'hFFFFFFF0;
    // rom_array[38564] = 32'hFFFFFFF0;
    // rom_array[38565] = 32'hFFFFFFF1;
    // rom_array[38566] = 32'hFFFFFFF1;
    // rom_array[38567] = 32'hFFFFFFF1;
    // rom_array[38568] = 32'hFFFFFFF1;
    // rom_array[38569] = 32'hFFFFFFF0;
    // rom_array[38570] = 32'hFFFFFFF0;
    // rom_array[38571] = 32'hFFFFFFF0;
    // rom_array[38572] = 32'hFFFFFFF0;
    // rom_array[38573] = 32'hFFFFFFF1;
    // rom_array[38574] = 32'hFFFFFFF1;
    // rom_array[38575] = 32'hFFFFFFF1;
    // rom_array[38576] = 32'hFFFFFFF1;
    // rom_array[38577] = 32'hFFFFFFF0;
    // rom_array[38578] = 32'hFFFFFFF0;
    // rom_array[38579] = 32'hFFFFFFF0;
    // rom_array[38580] = 32'hFFFFFFF0;
    // rom_array[38581] = 32'hFFFFFFF1;
    // rom_array[38582] = 32'hFFFFFFF1;
    // rom_array[38583] = 32'hFFFFFFF1;
    // rom_array[38584] = 32'hFFFFFFF1;
    // rom_array[38585] = 32'hFFFFFFF0;
    // rom_array[38586] = 32'hFFFFFFF0;
    // rom_array[38587] = 32'hFFFFFFF0;
    // rom_array[38588] = 32'hFFFFFFF0;
    // rom_array[38589] = 32'hFFFFFFF1;
    // rom_array[38590] = 32'hFFFFFFF1;
    // rom_array[38591] = 32'hFFFFFFF1;
    // rom_array[38592] = 32'hFFFFFFF1;
    // rom_array[38593] = 32'hFFFFFFF0;
    // rom_array[38594] = 32'hFFFFFFF0;
    // rom_array[38595] = 32'hFFFFFFF0;
    // rom_array[38596] = 32'hFFFFFFF0;
    // rom_array[38597] = 32'hFFFFFFF1;
    // rom_array[38598] = 32'hFFFFFFF1;
    // rom_array[38599] = 32'hFFFFFFF1;
    // rom_array[38600] = 32'hFFFFFFF1;
    // rom_array[38601] = 32'hFFFFFFF0;
    // rom_array[38602] = 32'hFFFFFFF0;
    // rom_array[38603] = 32'hFFFFFFF0;
    // rom_array[38604] = 32'hFFFFFFF0;
    // rom_array[38605] = 32'hFFFFFFF1;
    // rom_array[38606] = 32'hFFFFFFF1;
    // rom_array[38607] = 32'hFFFFFFF1;
    // rom_array[38608] = 32'hFFFFFFF1;
    // rom_array[38609] = 32'hFFFFFFF0;
    // rom_array[38610] = 32'hFFFFFFF0;
    // rom_array[38611] = 32'hFFFFFFF0;
    // rom_array[38612] = 32'hFFFFFFF0;
    // rom_array[38613] = 32'hFFFFFFF1;
    // rom_array[38614] = 32'hFFFFFFF1;
    // rom_array[38615] = 32'hFFFFFFF1;
    // rom_array[38616] = 32'hFFFFFFF1;
    // rom_array[38617] = 32'hFFFFFFF0;
    // rom_array[38618] = 32'hFFFFFFF0;
    // rom_array[38619] = 32'hFFFFFFF0;
    // rom_array[38620] = 32'hFFFFFFF0;
    // rom_array[38621] = 32'hFFFFFFF1;
    // rom_array[38622] = 32'hFFFFFFF1;
    // rom_array[38623] = 32'hFFFFFFF1;
    // rom_array[38624] = 32'hFFFFFFF1;
    // rom_array[38625] = 32'hFFFFFFF0;
    // rom_array[38626] = 32'hFFFFFFF0;
    // rom_array[38627] = 32'hFFFFFFF0;
    // rom_array[38628] = 32'hFFFFFFF0;
    // rom_array[38629] = 32'hFFFFFFF1;
    // rom_array[38630] = 32'hFFFFFFF1;
    // rom_array[38631] = 32'hFFFFFFF1;
    // rom_array[38632] = 32'hFFFFFFF1;
    // rom_array[38633] = 32'hFFFFFFF0;
    // rom_array[38634] = 32'hFFFFFFF0;
    // rom_array[38635] = 32'hFFFFFFF0;
    // rom_array[38636] = 32'hFFFFFFF0;
    // rom_array[38637] = 32'hFFFFFFF1;
    // rom_array[38638] = 32'hFFFFFFF1;
    // rom_array[38639] = 32'hFFFFFFF1;
    // rom_array[38640] = 32'hFFFFFFF1;
    // rom_array[38641] = 32'hFFFFFFF0;
    // rom_array[38642] = 32'hFFFFFFF0;
    // rom_array[38643] = 32'hFFFFFFF0;
    // rom_array[38644] = 32'hFFFFFFF0;
    // rom_array[38645] = 32'hFFFFFFF1;
    // rom_array[38646] = 32'hFFFFFFF1;
    // rom_array[38647] = 32'hFFFFFFF1;
    // rom_array[38648] = 32'hFFFFFFF1;
    // rom_array[38649] = 32'hFFFFFFF0;
    // rom_array[38650] = 32'hFFFFFFF0;
    // rom_array[38651] = 32'hFFFFFFF0;
    // rom_array[38652] = 32'hFFFFFFF0;
    // rom_array[38653] = 32'hFFFFFFF1;
    // rom_array[38654] = 32'hFFFFFFF1;
    // rom_array[38655] = 32'hFFFFFFF1;
    // rom_array[38656] = 32'hFFFFFFF1;
    // rom_array[38657] = 32'hFFFFFFF0;
    // rom_array[38658] = 32'hFFFFFFF0;
    // rom_array[38659] = 32'hFFFFFFF0;
    // rom_array[38660] = 32'hFFFFFFF0;
    // rom_array[38661] = 32'hFFFFFFF1;
    // rom_array[38662] = 32'hFFFFFFF1;
    // rom_array[38663] = 32'hFFFFFFF1;
    // rom_array[38664] = 32'hFFFFFFF1;
    // rom_array[38665] = 32'hFFFFFFF0;
    // rom_array[38666] = 32'hFFFFFFF0;
    // rom_array[38667] = 32'hFFFFFFF1;
    // rom_array[38668] = 32'hFFFFFFF1;
    // rom_array[38669] = 32'hFFFFFFF0;
    // rom_array[38670] = 32'hFFFFFFF0;
    // rom_array[38671] = 32'hFFFFFFF1;
    // rom_array[38672] = 32'hFFFFFFF1;
    // rom_array[38673] = 32'hFFFFFFF0;
    // rom_array[38674] = 32'hFFFFFFF0;
    // rom_array[38675] = 32'hFFFFFFF1;
    // rom_array[38676] = 32'hFFFFFFF1;
    // rom_array[38677] = 32'hFFFFFFF0;
    // rom_array[38678] = 32'hFFFFFFF0;
    // rom_array[38679] = 32'hFFFFFFF1;
    // rom_array[38680] = 32'hFFFFFFF1;
    // rom_array[38681] = 32'hFFFFFFF1;
    // rom_array[38682] = 32'hFFFFFFF1;
    // rom_array[38683] = 32'hFFFFFFF1;
    // rom_array[38684] = 32'hFFFFFFF1;
    // rom_array[38685] = 32'hFFFFFFF1;
    // rom_array[38686] = 32'hFFFFFFF1;
    // rom_array[38687] = 32'hFFFFFFF1;
    // rom_array[38688] = 32'hFFFFFFF1;
    // rom_array[38689] = 32'hFFFFFFF1;
    // rom_array[38690] = 32'hFFFFFFF1;
    // rom_array[38691] = 32'hFFFFFFF1;
    // rom_array[38692] = 32'hFFFFFFF1;
    // rom_array[38693] = 32'hFFFFFFF1;
    // rom_array[38694] = 32'hFFFFFFF1;
    // rom_array[38695] = 32'hFFFFFFF1;
    // rom_array[38696] = 32'hFFFFFFF1;
    // rom_array[38697] = 32'hFFFFFFF0;
    // rom_array[38698] = 32'hFFFFFFF0;
    // rom_array[38699] = 32'hFFFFFFF1;
    // rom_array[38700] = 32'hFFFFFFF1;
    // rom_array[38701] = 32'hFFFFFFF0;
    // rom_array[38702] = 32'hFFFFFFF0;
    // rom_array[38703] = 32'hFFFFFFF1;
    // rom_array[38704] = 32'hFFFFFFF1;
    // rom_array[38705] = 32'hFFFFFFF0;
    // rom_array[38706] = 32'hFFFFFFF0;
    // rom_array[38707] = 32'hFFFFFFF1;
    // rom_array[38708] = 32'hFFFFFFF1;
    // rom_array[38709] = 32'hFFFFFFF0;
    // rom_array[38710] = 32'hFFFFFFF0;
    // rom_array[38711] = 32'hFFFFFFF1;
    // rom_array[38712] = 32'hFFFFFFF1;
    // rom_array[38713] = 32'hFFFFFFF1;
    // rom_array[38714] = 32'hFFFFFFF1;
    // rom_array[38715] = 32'hFFFFFFF1;
    // rom_array[38716] = 32'hFFFFFFF1;
    // rom_array[38717] = 32'hFFFFFFF1;
    // rom_array[38718] = 32'hFFFFFFF1;
    // rom_array[38719] = 32'hFFFFFFF1;
    // rom_array[38720] = 32'hFFFFFFF1;
    // rom_array[38721] = 32'hFFFFFFF1;
    // rom_array[38722] = 32'hFFFFFFF1;
    // rom_array[38723] = 32'hFFFFFFF1;
    // rom_array[38724] = 32'hFFFFFFF1;
    // rom_array[38725] = 32'hFFFFFFF1;
    // rom_array[38726] = 32'hFFFFFFF1;
    // rom_array[38727] = 32'hFFFFFFF1;
    // rom_array[38728] = 32'hFFFFFFF1;
    // rom_array[38729] = 32'hFFFFFFF1;
    // rom_array[38730] = 32'hFFFFFFF1;
    // rom_array[38731] = 32'hFFFFFFF1;
    // rom_array[38732] = 32'hFFFFFFF1;
    // rom_array[38733] = 32'hFFFFFFF1;
    // rom_array[38734] = 32'hFFFFFFF1;
    // rom_array[38735] = 32'hFFFFFFF1;
    // rom_array[38736] = 32'hFFFFFFF1;
    // rom_array[38737] = 32'hFFFFFFF1;
    // rom_array[38738] = 32'hFFFFFFF1;
    // rom_array[38739] = 32'hFFFFFFF1;
    // rom_array[38740] = 32'hFFFFFFF1;
    // rom_array[38741] = 32'hFFFFFFF1;
    // rom_array[38742] = 32'hFFFFFFF1;
    // rom_array[38743] = 32'hFFFFFFF1;
    // rom_array[38744] = 32'hFFFFFFF1;
    // rom_array[38745] = 32'hFFFFFFF0;
    // rom_array[38746] = 32'hFFFFFFF0;
    // rom_array[38747] = 32'hFFFFFFF1;
    // rom_array[38748] = 32'hFFFFFFF1;
    // rom_array[38749] = 32'hFFFFFFF0;
    // rom_array[38750] = 32'hFFFFFFF0;
    // rom_array[38751] = 32'hFFFFFFF1;
    // rom_array[38752] = 32'hFFFFFFF1;
    // rom_array[38753] = 32'hFFFFFFF0;
    // rom_array[38754] = 32'hFFFFFFF0;
    // rom_array[38755] = 32'hFFFFFFF1;
    // rom_array[38756] = 32'hFFFFFFF1;
    // rom_array[38757] = 32'hFFFFFFF0;
    // rom_array[38758] = 32'hFFFFFFF0;
    // rom_array[38759] = 32'hFFFFFFF1;
    // rom_array[38760] = 32'hFFFFFFF1;
    // rom_array[38761] = 32'hFFFFFFF0;
    // rom_array[38762] = 32'hFFFFFFF0;
    // rom_array[38763] = 32'hFFFFFFF1;
    // rom_array[38764] = 32'hFFFFFFF1;
    // rom_array[38765] = 32'hFFFFFFF0;
    // rom_array[38766] = 32'hFFFFFFF0;
    // rom_array[38767] = 32'hFFFFFFF1;
    // rom_array[38768] = 32'hFFFFFFF1;
    // rom_array[38769] = 32'hFFFFFFF0;
    // rom_array[38770] = 32'hFFFFFFF0;
    // rom_array[38771] = 32'hFFFFFFF1;
    // rom_array[38772] = 32'hFFFFFFF1;
    // rom_array[38773] = 32'hFFFFFFF0;
    // rom_array[38774] = 32'hFFFFFFF0;
    // rom_array[38775] = 32'hFFFFFFF1;
    // rom_array[38776] = 32'hFFFFFFF1;
    // rom_array[38777] = 32'hFFFFFFF0;
    // rom_array[38778] = 32'hFFFFFFF0;
    // rom_array[38779] = 32'hFFFFFFF1;
    // rom_array[38780] = 32'hFFFFFFF1;
    // rom_array[38781] = 32'hFFFFFFF0;
    // rom_array[38782] = 32'hFFFFFFF0;
    // rom_array[38783] = 32'hFFFFFFF1;
    // rom_array[38784] = 32'hFFFFFFF1;
    // rom_array[38785] = 32'hFFFFFFF0;
    // rom_array[38786] = 32'hFFFFFFF0;
    // rom_array[38787] = 32'hFFFFFFF1;
    // rom_array[38788] = 32'hFFFFFFF1;
    // rom_array[38789] = 32'hFFFFFFF0;
    // rom_array[38790] = 32'hFFFFFFF0;
    // rom_array[38791] = 32'hFFFFFFF1;
    // rom_array[38792] = 32'hFFFFFFF1;
    // rom_array[38793] = 32'hFFFFFFF0;
    // rom_array[38794] = 32'hFFFFFFF0;
    // rom_array[38795] = 32'hFFFFFFF1;
    // rom_array[38796] = 32'hFFFFFFF1;
    // rom_array[38797] = 32'hFFFFFFF0;
    // rom_array[38798] = 32'hFFFFFFF0;
    // rom_array[38799] = 32'hFFFFFFF1;
    // rom_array[38800] = 32'hFFFFFFF1;
    // rom_array[38801] = 32'hFFFFFFF0;
    // rom_array[38802] = 32'hFFFFFFF0;
    // rom_array[38803] = 32'hFFFFFFF1;
    // rom_array[38804] = 32'hFFFFFFF1;
    // rom_array[38805] = 32'hFFFFFFF0;
    // rom_array[38806] = 32'hFFFFFFF0;
    // rom_array[38807] = 32'hFFFFFFF1;
    // rom_array[38808] = 32'hFFFFFFF1;
    // rom_array[38809] = 32'hFFFFFFF0;
    // rom_array[38810] = 32'hFFFFFFF0;
    // rom_array[38811] = 32'hFFFFFFF1;
    // rom_array[38812] = 32'hFFFFFFF1;
    // rom_array[38813] = 32'hFFFFFFF0;
    // rom_array[38814] = 32'hFFFFFFF0;
    // rom_array[38815] = 32'hFFFFFFF1;
    // rom_array[38816] = 32'hFFFFFFF1;
    // rom_array[38817] = 32'hFFFFFFF0;
    // rom_array[38818] = 32'hFFFFFFF0;
    // rom_array[38819] = 32'hFFFFFFF1;
    // rom_array[38820] = 32'hFFFFFFF1;
    // rom_array[38821] = 32'hFFFFFFF0;
    // rom_array[38822] = 32'hFFFFFFF0;
    // rom_array[38823] = 32'hFFFFFFF1;
    // rom_array[38824] = 32'hFFFFFFF1;
    // rom_array[38825] = 32'hFFFFFFF0;
    // rom_array[38826] = 32'hFFFFFFF0;
    // rom_array[38827] = 32'hFFFFFFF1;
    // rom_array[38828] = 32'hFFFFFFF1;
    // rom_array[38829] = 32'hFFFFFFF0;
    // rom_array[38830] = 32'hFFFFFFF0;
    // rom_array[38831] = 32'hFFFFFFF1;
    // rom_array[38832] = 32'hFFFFFFF1;
    // rom_array[38833] = 32'hFFFFFFF0;
    // rom_array[38834] = 32'hFFFFFFF0;
    // rom_array[38835] = 32'hFFFFFFF1;
    // rom_array[38836] = 32'hFFFFFFF1;
    // rom_array[38837] = 32'hFFFFFFF0;
    // rom_array[38838] = 32'hFFFFFFF0;
    // rom_array[38839] = 32'hFFFFFFF1;
    // rom_array[38840] = 32'hFFFFFFF1;
    // rom_array[38841] = 32'hFFFFFFF1;
    // rom_array[38842] = 32'hFFFFFFF1;
    // rom_array[38843] = 32'hFFFFFFF1;
    // rom_array[38844] = 32'hFFFFFFF1;
    // rom_array[38845] = 32'hFFFFFFF1;
    // rom_array[38846] = 32'hFFFFFFF1;
    // rom_array[38847] = 32'hFFFFFFF1;
    // rom_array[38848] = 32'hFFFFFFF1;
    // rom_array[38849] = 32'hFFFFFFF1;
    // rom_array[38850] = 32'hFFFFFFF1;
    // rom_array[38851] = 32'hFFFFFFF1;
    // rom_array[38852] = 32'hFFFFFFF1;
    // rom_array[38853] = 32'hFFFFFFF1;
    // rom_array[38854] = 32'hFFFFFFF1;
    // rom_array[38855] = 32'hFFFFFFF1;
    // rom_array[38856] = 32'hFFFFFFF1;
    // rom_array[38857] = 32'hFFFFFFF1;
    // rom_array[38858] = 32'hFFFFFFF1;
    // rom_array[38859] = 32'hFFFFFFF1;
    // rom_array[38860] = 32'hFFFFFFF1;
    // rom_array[38861] = 32'hFFFFFFF0;
    // rom_array[38862] = 32'hFFFFFFF0;
    // rom_array[38863] = 32'hFFFFFFF0;
    // rom_array[38864] = 32'hFFFFFFF0;
    // rom_array[38865] = 32'hFFFFFFF1;
    // rom_array[38866] = 32'hFFFFFFF1;
    // rom_array[38867] = 32'hFFFFFFF1;
    // rom_array[38868] = 32'hFFFFFFF1;
    // rom_array[38869] = 32'hFFFFFFF0;
    // rom_array[38870] = 32'hFFFFFFF0;
    // rom_array[38871] = 32'hFFFFFFF0;
    // rom_array[38872] = 32'hFFFFFFF0;
    // rom_array[38873] = 32'hFFFFFFF1;
    // rom_array[38874] = 32'hFFFFFFF1;
    // rom_array[38875] = 32'hFFFFFFF1;
    // rom_array[38876] = 32'hFFFFFFF1;
    // rom_array[38877] = 32'hFFFFFFF1;
    // rom_array[38878] = 32'hFFFFFFF1;
    // rom_array[38879] = 32'hFFFFFFF1;
    // rom_array[38880] = 32'hFFFFFFF1;
    // rom_array[38881] = 32'hFFFFFFF1;
    // rom_array[38882] = 32'hFFFFFFF1;
    // rom_array[38883] = 32'hFFFFFFF1;
    // rom_array[38884] = 32'hFFFFFFF1;
    // rom_array[38885] = 32'hFFFFFFF1;
    // rom_array[38886] = 32'hFFFFFFF1;
    // rom_array[38887] = 32'hFFFFFFF1;
    // rom_array[38888] = 32'hFFFFFFF1;
    // rom_array[38889] = 32'hFFFFFFF1;
    // rom_array[38890] = 32'hFFFFFFF1;
    // rom_array[38891] = 32'hFFFFFFF1;
    // rom_array[38892] = 32'hFFFFFFF1;
    // rom_array[38893] = 32'hFFFFFFF0;
    // rom_array[38894] = 32'hFFFFFFF0;
    // rom_array[38895] = 32'hFFFFFFF0;
    // rom_array[38896] = 32'hFFFFFFF0;
    // rom_array[38897] = 32'hFFFFFFF1;
    // rom_array[38898] = 32'hFFFFFFF1;
    // rom_array[38899] = 32'hFFFFFFF1;
    // rom_array[38900] = 32'hFFFFFFF1;
    // rom_array[38901] = 32'hFFFFFFF0;
    // rom_array[38902] = 32'hFFFFFFF0;
    // rom_array[38903] = 32'hFFFFFFF0;
    // rom_array[38904] = 32'hFFFFFFF0;
    // rom_array[38905] = 32'hFFFFFFF1;
    // rom_array[38906] = 32'hFFFFFFF1;
    // rom_array[38907] = 32'hFFFFFFF1;
    // rom_array[38908] = 32'hFFFFFFF1;
    // rom_array[38909] = 32'hFFFFFFF0;
    // rom_array[38910] = 32'hFFFFFFF0;
    // rom_array[38911] = 32'hFFFFFFF0;
    // rom_array[38912] = 32'hFFFFFFF0;
    // rom_array[38913] = 32'hFFFFFFF1;
    // rom_array[38914] = 32'hFFFFFFF1;
    // rom_array[38915] = 32'hFFFFFFF1;
    // rom_array[38916] = 32'hFFFFFFF1;
    // rom_array[38917] = 32'hFFFFFFF0;
    // rom_array[38918] = 32'hFFFFFFF0;
    // rom_array[38919] = 32'hFFFFFFF0;
    // rom_array[38920] = 32'hFFFFFFF0;
    // rom_array[38921] = 32'hFFFFFFF1;
    // rom_array[38922] = 32'hFFFFFFF1;
    // rom_array[38923] = 32'hFFFFFFF1;
    // rom_array[38924] = 32'hFFFFFFF1;
    // rom_array[38925] = 32'hFFFFFFF1;
    // rom_array[38926] = 32'hFFFFFFF1;
    // rom_array[38927] = 32'hFFFFFFF1;
    // rom_array[38928] = 32'hFFFFFFF1;
    // rom_array[38929] = 32'hFFFFFFF1;
    // rom_array[38930] = 32'hFFFFFFF1;
    // rom_array[38931] = 32'hFFFFFFF1;
    // rom_array[38932] = 32'hFFFFFFF1;
    // rom_array[38933] = 32'hFFFFFFF1;
    // rom_array[38934] = 32'hFFFFFFF1;
    // rom_array[38935] = 32'hFFFFFFF1;
    // rom_array[38936] = 32'hFFFFFFF1;
    // rom_array[38937] = 32'hFFFFFFF1;
    // rom_array[38938] = 32'hFFFFFFF1;
    // rom_array[38939] = 32'hFFFFFFF1;
    // rom_array[38940] = 32'hFFFFFFF1;
    // rom_array[38941] = 32'hFFFFFFF1;
    // rom_array[38942] = 32'hFFFFFFF1;
    // rom_array[38943] = 32'hFFFFFFF1;
    // rom_array[38944] = 32'hFFFFFFF1;
    // rom_array[38945] = 32'hFFFFFFF1;
    // rom_array[38946] = 32'hFFFFFFF1;
    // rom_array[38947] = 32'hFFFFFFF1;
    // rom_array[38948] = 32'hFFFFFFF1;
    // rom_array[38949] = 32'hFFFFFFF1;
    // rom_array[38950] = 32'hFFFFFFF1;
    // rom_array[38951] = 32'hFFFFFFF1;
    // rom_array[38952] = 32'hFFFFFFF1;
    // rom_array[38953] = 32'hFFFFFFF1;
    // rom_array[38954] = 32'hFFFFFFF1;
    // rom_array[38955] = 32'hFFFFFFF1;
    // rom_array[38956] = 32'hFFFFFFF1;
    // rom_array[38957] = 32'hFFFFFFF0;
    // rom_array[38958] = 32'hFFFFFFF0;
    // rom_array[38959] = 32'hFFFFFFF0;
    // rom_array[38960] = 32'hFFFFFFF0;
    // rom_array[38961] = 32'hFFFFFFF1;
    // rom_array[38962] = 32'hFFFFFFF1;
    // rom_array[38963] = 32'hFFFFFFF1;
    // rom_array[38964] = 32'hFFFFFFF1;
    // rom_array[38965] = 32'hFFFFFFF0;
    // rom_array[38966] = 32'hFFFFFFF0;
    // rom_array[38967] = 32'hFFFFFFF0;
    // rom_array[38968] = 32'hFFFFFFF0;
    // rom_array[38969] = 32'hFFFFFFF1;
    // rom_array[38970] = 32'hFFFFFFF1;
    // rom_array[38971] = 32'hFFFFFFF1;
    // rom_array[38972] = 32'hFFFFFFF1;
    // rom_array[38973] = 32'hFFFFFFF0;
    // rom_array[38974] = 32'hFFFFFFF0;
    // rom_array[38975] = 32'hFFFFFFF0;
    // rom_array[38976] = 32'hFFFFFFF0;
    // rom_array[38977] = 32'hFFFFFFF1;
    // rom_array[38978] = 32'hFFFFFFF1;
    // rom_array[38979] = 32'hFFFFFFF1;
    // rom_array[38980] = 32'hFFFFFFF1;
    // rom_array[38981] = 32'hFFFFFFF0;
    // rom_array[38982] = 32'hFFFFFFF0;
    // rom_array[38983] = 32'hFFFFFFF0;
    // rom_array[38984] = 32'hFFFFFFF0;
    // rom_array[38985] = 32'hFFFFFFF1;
    // rom_array[38986] = 32'hFFFFFFF1;
    // rom_array[38987] = 32'hFFFFFFF1;
    // rom_array[38988] = 32'hFFFFFFF1;
    // rom_array[38989] = 32'hFFFFFFF0;
    // rom_array[38990] = 32'hFFFFFFF0;
    // rom_array[38991] = 32'hFFFFFFF0;
    // rom_array[38992] = 32'hFFFFFFF0;
    // rom_array[38993] = 32'hFFFFFFF1;
    // rom_array[38994] = 32'hFFFFFFF1;
    // rom_array[38995] = 32'hFFFFFFF1;
    // rom_array[38996] = 32'hFFFFFFF1;
    // rom_array[38997] = 32'hFFFFFFF0;
    // rom_array[38998] = 32'hFFFFFFF0;
    // rom_array[38999] = 32'hFFFFFFF0;
    // rom_array[39000] = 32'hFFFFFFF0;
    // rom_array[39001] = 32'hFFFFFFF1;
    // rom_array[39002] = 32'hFFFFFFF1;
    // rom_array[39003] = 32'hFFFFFFF1;
    // rom_array[39004] = 32'hFFFFFFF1;
    // rom_array[39005] = 32'hFFFFFFF0;
    // rom_array[39006] = 32'hFFFFFFF0;
    // rom_array[39007] = 32'hFFFFFFF0;
    // rom_array[39008] = 32'hFFFFFFF0;
    // rom_array[39009] = 32'hFFFFFFF1;
    // rom_array[39010] = 32'hFFFFFFF1;
    // rom_array[39011] = 32'hFFFFFFF1;
    // rom_array[39012] = 32'hFFFFFFF1;
    // rom_array[39013] = 32'hFFFFFFF0;
    // rom_array[39014] = 32'hFFFFFFF0;
    // rom_array[39015] = 32'hFFFFFFF0;
    // rom_array[39016] = 32'hFFFFFFF0;
    // rom_array[39017] = 32'hFFFFFFF1;
    // rom_array[39018] = 32'hFFFFFFF1;
    // rom_array[39019] = 32'hFFFFFFF1;
    // rom_array[39020] = 32'hFFFFFFF1;
    // rom_array[39021] = 32'hFFFFFFF1;
    // rom_array[39022] = 32'hFFFFFFF1;
    // rom_array[39023] = 32'hFFFFFFF1;
    // rom_array[39024] = 32'hFFFFFFF1;
    // rom_array[39025] = 32'hFFFFFFF1;
    // rom_array[39026] = 32'hFFFFFFF1;
    // rom_array[39027] = 32'hFFFFFFF1;
    // rom_array[39028] = 32'hFFFFFFF1;
    // rom_array[39029] = 32'hFFFFFFF1;
    // rom_array[39030] = 32'hFFFFFFF1;
    // rom_array[39031] = 32'hFFFFFFF1;
    // rom_array[39032] = 32'hFFFFFFF1;
    // rom_array[39033] = 32'hFFFFFFF1;
    // rom_array[39034] = 32'hFFFFFFF1;
    // rom_array[39035] = 32'hFFFFFFF1;
    // rom_array[39036] = 32'hFFFFFFF1;
    // rom_array[39037] = 32'hFFFFFFF1;
    // rom_array[39038] = 32'hFFFFFFF1;
    // rom_array[39039] = 32'hFFFFFFF1;
    // rom_array[39040] = 32'hFFFFFFF1;
    // rom_array[39041] = 32'hFFFFFFF1;
    // rom_array[39042] = 32'hFFFFFFF1;
    // rom_array[39043] = 32'hFFFFFFF1;
    // rom_array[39044] = 32'hFFFFFFF1;
    // rom_array[39045] = 32'hFFFFFFF1;
    // rom_array[39046] = 32'hFFFFFFF1;
    // rom_array[39047] = 32'hFFFFFFF1;
    // rom_array[39048] = 32'hFFFFFFF1;
    // rom_array[39049] = 32'hFFFFFFF1;
    // rom_array[39050] = 32'hFFFFFFF1;
    // rom_array[39051] = 32'hFFFFFFF1;
    // rom_array[39052] = 32'hFFFFFFF1;
    // rom_array[39053] = 32'hFFFFFFF1;
    // rom_array[39054] = 32'hFFFFFFF1;
    // rom_array[39055] = 32'hFFFFFFF1;
    // rom_array[39056] = 32'hFFFFFFF1;
    // rom_array[39057] = 32'hFFFFFFF1;
    // rom_array[39058] = 32'hFFFFFFF1;
    // rom_array[39059] = 32'hFFFFFFF1;
    // rom_array[39060] = 32'hFFFFFFF1;
    // rom_array[39061] = 32'hFFFFFFF1;
    // rom_array[39062] = 32'hFFFFFFF1;
    // rom_array[39063] = 32'hFFFFFFF1;
    // rom_array[39064] = 32'hFFFFFFF1;
    // rom_array[39065] = 32'hFFFFFFF1;
    // rom_array[39066] = 32'hFFFFFFF1;
    // rom_array[39067] = 32'hFFFFFFF1;
    // rom_array[39068] = 32'hFFFFFFF1;
    // rom_array[39069] = 32'hFFFFFFF1;
    // rom_array[39070] = 32'hFFFFFFF1;
    // rom_array[39071] = 32'hFFFFFFF1;
    // rom_array[39072] = 32'hFFFFFFF1;
    // rom_array[39073] = 32'hFFFFFFF1;
    // rom_array[39074] = 32'hFFFFFFF1;
    // rom_array[39075] = 32'hFFFFFFF1;
    // rom_array[39076] = 32'hFFFFFFF1;
    // rom_array[39077] = 32'hFFFFFFF1;
    // rom_array[39078] = 32'hFFFFFFF1;
    // rom_array[39079] = 32'hFFFFFFF1;
    // rom_array[39080] = 32'hFFFFFFF1;
    // rom_array[39081] = 32'hFFFFFFF0;
    // rom_array[39082] = 32'hFFFFFFF0;
    // rom_array[39083] = 32'hFFFFFFF1;
    // rom_array[39084] = 32'hFFFFFFF1;
    // rom_array[39085] = 32'hFFFFFFF0;
    // rom_array[39086] = 32'hFFFFFFF0;
    // rom_array[39087] = 32'hFFFFFFF1;
    // rom_array[39088] = 32'hFFFFFFF1;
    // rom_array[39089] = 32'hFFFFFFF0;
    // rom_array[39090] = 32'hFFFFFFF0;
    // rom_array[39091] = 32'hFFFFFFF1;
    // rom_array[39092] = 32'hFFFFFFF1;
    // rom_array[39093] = 32'hFFFFFFF0;
    // rom_array[39094] = 32'hFFFFFFF0;
    // rom_array[39095] = 32'hFFFFFFF1;
    // rom_array[39096] = 32'hFFFFFFF1;
    // rom_array[39097] = 32'hFFFFFFF0;
    // rom_array[39098] = 32'hFFFFFFF0;
    // rom_array[39099] = 32'hFFFFFFF1;
    // rom_array[39100] = 32'hFFFFFFF1;
    // rom_array[39101] = 32'hFFFFFFF0;
    // rom_array[39102] = 32'hFFFFFFF0;
    // rom_array[39103] = 32'hFFFFFFF1;
    // rom_array[39104] = 32'hFFFFFFF1;
    // rom_array[39105] = 32'hFFFFFFF0;
    // rom_array[39106] = 32'hFFFFFFF0;
    // rom_array[39107] = 32'hFFFFFFF1;
    // rom_array[39108] = 32'hFFFFFFF1;
    // rom_array[39109] = 32'hFFFFFFF0;
    // rom_array[39110] = 32'hFFFFFFF0;
    // rom_array[39111] = 32'hFFFFFFF1;
    // rom_array[39112] = 32'hFFFFFFF1;
    // rom_array[39113] = 32'hFFFFFFF0;
    // rom_array[39114] = 32'hFFFFFFF0;
    // rom_array[39115] = 32'hFFFFFFF1;
    // rom_array[39116] = 32'hFFFFFFF1;
    // rom_array[39117] = 32'hFFFFFFF0;
    // rom_array[39118] = 32'hFFFFFFF0;
    // rom_array[39119] = 32'hFFFFFFF0;
    // rom_array[39120] = 32'hFFFFFFF0;
    // rom_array[39121] = 32'hFFFFFFF0;
    // rom_array[39122] = 32'hFFFFFFF0;
    // rom_array[39123] = 32'hFFFFFFF1;
    // rom_array[39124] = 32'hFFFFFFF1;
    // rom_array[39125] = 32'hFFFFFFF0;
    // rom_array[39126] = 32'hFFFFFFF0;
    // rom_array[39127] = 32'hFFFFFFF0;
    // rom_array[39128] = 32'hFFFFFFF0;
    // rom_array[39129] = 32'hFFFFFFF1;
    // rom_array[39130] = 32'hFFFFFFF1;
    // rom_array[39131] = 32'hFFFFFFF1;
    // rom_array[39132] = 32'hFFFFFFF1;
    // rom_array[39133] = 32'hFFFFFFF0;
    // rom_array[39134] = 32'hFFFFFFF0;
    // rom_array[39135] = 32'hFFFFFFF0;
    // rom_array[39136] = 32'hFFFFFFF0;
    // rom_array[39137] = 32'hFFFFFFF1;
    // rom_array[39138] = 32'hFFFFFFF1;
    // rom_array[39139] = 32'hFFFFFFF1;
    // rom_array[39140] = 32'hFFFFFFF1;
    // rom_array[39141] = 32'hFFFFFFF0;
    // rom_array[39142] = 32'hFFFFFFF0;
    // rom_array[39143] = 32'hFFFFFFF0;
    // rom_array[39144] = 32'hFFFFFFF0;
    // rom_array[39145] = 32'hFFFFFFF1;
    // rom_array[39146] = 32'hFFFFFFF1;
    // rom_array[39147] = 32'hFFFFFFF1;
    // rom_array[39148] = 32'hFFFFFFF1;
    // rom_array[39149] = 32'hFFFFFFF0;
    // rom_array[39150] = 32'hFFFFFFF0;
    // rom_array[39151] = 32'hFFFFFFF0;
    // rom_array[39152] = 32'hFFFFFFF0;
    // rom_array[39153] = 32'hFFFFFFF1;
    // rom_array[39154] = 32'hFFFFFFF1;
    // rom_array[39155] = 32'hFFFFFFF1;
    // rom_array[39156] = 32'hFFFFFFF1;
    // rom_array[39157] = 32'hFFFFFFF0;
    // rom_array[39158] = 32'hFFFFFFF0;
    // rom_array[39159] = 32'hFFFFFFF0;
    // rom_array[39160] = 32'hFFFFFFF0;
    // rom_array[39161] = 32'hFFFFFFF1;
    // rom_array[39162] = 32'hFFFFFFF1;
    // rom_array[39163] = 32'hFFFFFFF1;
    // rom_array[39164] = 32'hFFFFFFF1;
    // rom_array[39165] = 32'hFFFFFFF0;
    // rom_array[39166] = 32'hFFFFFFF0;
    // rom_array[39167] = 32'hFFFFFFF0;
    // rom_array[39168] = 32'hFFFFFFF0;
    // rom_array[39169] = 32'hFFFFFFF1;
    // rom_array[39170] = 32'hFFFFFFF1;
    // rom_array[39171] = 32'hFFFFFFF1;
    // rom_array[39172] = 32'hFFFFFFF1;
    // rom_array[39173] = 32'hFFFFFFF0;
    // rom_array[39174] = 32'hFFFFFFF0;
    // rom_array[39175] = 32'hFFFFFFF0;
    // rom_array[39176] = 32'hFFFFFFF0;
    // rom_array[39177] = 32'hFFFFFFF1;
    // rom_array[39178] = 32'hFFFFFFF1;
    // rom_array[39179] = 32'hFFFFFFF1;
    // rom_array[39180] = 32'hFFFFFFF1;
    // rom_array[39181] = 32'hFFFFFFF1;
    // rom_array[39182] = 32'hFFFFFFF1;
    // rom_array[39183] = 32'hFFFFFFF1;
    // rom_array[39184] = 32'hFFFFFFF1;
    // rom_array[39185] = 32'hFFFFFFF1;
    // rom_array[39186] = 32'hFFFFFFF1;
    // rom_array[39187] = 32'hFFFFFFF1;
    // rom_array[39188] = 32'hFFFFFFF1;
    // rom_array[39189] = 32'hFFFFFFF1;
    // rom_array[39190] = 32'hFFFFFFF1;
    // rom_array[39191] = 32'hFFFFFFF1;
    // rom_array[39192] = 32'hFFFFFFF1;
    // rom_array[39193] = 32'hFFFFFFF1;
    // rom_array[39194] = 32'hFFFFFFF1;
    // rom_array[39195] = 32'hFFFFFFF1;
    // rom_array[39196] = 32'hFFFFFFF1;
    // rom_array[39197] = 32'hFFFFFFF1;
    // rom_array[39198] = 32'hFFFFFFF1;
    // rom_array[39199] = 32'hFFFFFFF1;
    // rom_array[39200] = 32'hFFFFFFF1;
    // rom_array[39201] = 32'hFFFFFFF1;
    // rom_array[39202] = 32'hFFFFFFF1;
    // rom_array[39203] = 32'hFFFFFFF1;
    // rom_array[39204] = 32'hFFFFFFF1;
    // rom_array[39205] = 32'hFFFFFFF1;
    // rom_array[39206] = 32'hFFFFFFF1;
    // rom_array[39207] = 32'hFFFFFFF1;
    // rom_array[39208] = 32'hFFFFFFF1;
    // rom_array[39209] = 32'hFFFFFFF1;
    // rom_array[39210] = 32'hFFFFFFF1;
    // rom_array[39211] = 32'hFFFFFFF1;
    // rom_array[39212] = 32'hFFFFFFF1;
    // rom_array[39213] = 32'hFFFFFFF0;
    // rom_array[39214] = 32'hFFFFFFF0;
    // rom_array[39215] = 32'hFFFFFFF0;
    // rom_array[39216] = 32'hFFFFFFF0;
    // rom_array[39217] = 32'hFFFFFFF1;
    // rom_array[39218] = 32'hFFFFFFF1;
    // rom_array[39219] = 32'hFFFFFFF1;
    // rom_array[39220] = 32'hFFFFFFF1;
    // rom_array[39221] = 32'hFFFFFFF0;
    // rom_array[39222] = 32'hFFFFFFF0;
    // rom_array[39223] = 32'hFFFFFFF0;
    // rom_array[39224] = 32'hFFFFFFF0;
    // rom_array[39225] = 32'hFFFFFFF1;
    // rom_array[39226] = 32'hFFFFFFF1;
    // rom_array[39227] = 32'hFFFFFFF1;
    // rom_array[39228] = 32'hFFFFFFF1;
    // rom_array[39229] = 32'hFFFFFFF0;
    // rom_array[39230] = 32'hFFFFFFF0;
    // rom_array[39231] = 32'hFFFFFFF0;
    // rom_array[39232] = 32'hFFFFFFF0;
    // rom_array[39233] = 32'hFFFFFFF1;
    // rom_array[39234] = 32'hFFFFFFF1;
    // rom_array[39235] = 32'hFFFFFFF1;
    // rom_array[39236] = 32'hFFFFFFF1;
    // rom_array[39237] = 32'hFFFFFFF0;
    // rom_array[39238] = 32'hFFFFFFF0;
    // rom_array[39239] = 32'hFFFFFFF0;
    // rom_array[39240] = 32'hFFFFFFF0;
    // rom_array[39241] = 32'hFFFFFFF1;
    // rom_array[39242] = 32'hFFFFFFF1;
    // rom_array[39243] = 32'hFFFFFFF1;
    // rom_array[39244] = 32'hFFFFFFF1;
    // rom_array[39245] = 32'hFFFFFFF0;
    // rom_array[39246] = 32'hFFFFFFF0;
    // rom_array[39247] = 32'hFFFFFFF0;
    // rom_array[39248] = 32'hFFFFFFF0;
    // rom_array[39249] = 32'hFFFFFFF1;
    // rom_array[39250] = 32'hFFFFFFF1;
    // rom_array[39251] = 32'hFFFFFFF1;
    // rom_array[39252] = 32'hFFFFFFF1;
    // rom_array[39253] = 32'hFFFFFFF0;
    // rom_array[39254] = 32'hFFFFFFF0;
    // rom_array[39255] = 32'hFFFFFFF0;
    // rom_array[39256] = 32'hFFFFFFF0;
    // rom_array[39257] = 32'hFFFFFFF0;
    // rom_array[39258] = 32'hFFFFFFF0;
    // rom_array[39259] = 32'hFFFFFFF1;
    // rom_array[39260] = 32'hFFFFFFF1;
    // rom_array[39261] = 32'hFFFFFFF0;
    // rom_array[39262] = 32'hFFFFFFF0;
    // rom_array[39263] = 32'hFFFFFFF0;
    // rom_array[39264] = 32'hFFFFFFF0;
    // rom_array[39265] = 32'hFFFFFFF0;
    // rom_array[39266] = 32'hFFFFFFF0;
    // rom_array[39267] = 32'hFFFFFFF1;
    // rom_array[39268] = 32'hFFFFFFF1;
    // rom_array[39269] = 32'hFFFFFFF0;
    // rom_array[39270] = 32'hFFFFFFF0;
    // rom_array[39271] = 32'hFFFFFFF0;
    // rom_array[39272] = 32'hFFFFFFF0;
    // rom_array[39273] = 32'hFFFFFFF1;
    // rom_array[39274] = 32'hFFFFFFF1;
    // rom_array[39275] = 32'hFFFFFFF1;
    // rom_array[39276] = 32'hFFFFFFF1;
    // rom_array[39277] = 32'hFFFFFFF0;
    // rom_array[39278] = 32'hFFFFFFF0;
    // rom_array[39279] = 32'hFFFFFFF0;
    // rom_array[39280] = 32'hFFFFFFF0;
    // rom_array[39281] = 32'hFFFFFFF1;
    // rom_array[39282] = 32'hFFFFFFF1;
    // rom_array[39283] = 32'hFFFFFFF1;
    // rom_array[39284] = 32'hFFFFFFF1;
    // rom_array[39285] = 32'hFFFFFFF0;
    // rom_array[39286] = 32'hFFFFFFF0;
    // rom_array[39287] = 32'hFFFFFFF0;
    // rom_array[39288] = 32'hFFFFFFF0;
    // rom_array[39289] = 32'hFFFFFFF1;
    // rom_array[39290] = 32'hFFFFFFF1;
    // rom_array[39291] = 32'hFFFFFFF1;
    // rom_array[39292] = 32'hFFFFFFF1;
    // rom_array[39293] = 32'hFFFFFFF0;
    // rom_array[39294] = 32'hFFFFFFF0;
    // rom_array[39295] = 32'hFFFFFFF0;
    // rom_array[39296] = 32'hFFFFFFF0;
    // rom_array[39297] = 32'hFFFFFFF1;
    // rom_array[39298] = 32'hFFFFFFF1;
    // rom_array[39299] = 32'hFFFFFFF1;
    // rom_array[39300] = 32'hFFFFFFF1;
    // rom_array[39301] = 32'hFFFFFFF0;
    // rom_array[39302] = 32'hFFFFFFF0;
    // rom_array[39303] = 32'hFFFFFFF0;
    // rom_array[39304] = 32'hFFFFFFF0;
    // rom_array[39305] = 32'hFFFFFFF1;
    // rom_array[39306] = 32'hFFFFFFF1;
    // rom_array[39307] = 32'hFFFFFFF1;
    // rom_array[39308] = 32'hFFFFFFF1;
    // rom_array[39309] = 32'hFFFFFFF0;
    // rom_array[39310] = 32'hFFFFFFF0;
    // rom_array[39311] = 32'hFFFFFFF0;
    // rom_array[39312] = 32'hFFFFFFF0;
    // rom_array[39313] = 32'hFFFFFFF1;
    // rom_array[39314] = 32'hFFFFFFF1;
    // rom_array[39315] = 32'hFFFFFFF1;
    // rom_array[39316] = 32'hFFFFFFF1;
    // rom_array[39317] = 32'hFFFFFFF0;
    // rom_array[39318] = 32'hFFFFFFF0;
    // rom_array[39319] = 32'hFFFFFFF0;
    // rom_array[39320] = 32'hFFFFFFF0;
    // rom_array[39321] = 32'hFFFFFFF1;
    // rom_array[39322] = 32'hFFFFFFF1;
    // rom_array[39323] = 32'hFFFFFFF1;
    // rom_array[39324] = 32'hFFFFFFF1;
    // rom_array[39325] = 32'hFFFFFFF0;
    // rom_array[39326] = 32'hFFFFFFF0;
    // rom_array[39327] = 32'hFFFFFFF0;
    // rom_array[39328] = 32'hFFFFFFF0;
    // rom_array[39329] = 32'hFFFFFFF1;
    // rom_array[39330] = 32'hFFFFFFF1;
    // rom_array[39331] = 32'hFFFFFFF1;
    // rom_array[39332] = 32'hFFFFFFF1;
    // rom_array[39333] = 32'hFFFFFFF0;
    // rom_array[39334] = 32'hFFFFFFF0;
    // rom_array[39335] = 32'hFFFFFFF0;
    // rom_array[39336] = 32'hFFFFFFF0;
    // rom_array[39337] = 32'hFFFFFFF0;
    // rom_array[39338] = 32'hFFFFFFF0;
    // rom_array[39339] = 32'hFFFFFFF0;
    // rom_array[39340] = 32'hFFFFFFF0;
    // rom_array[39341] = 32'hFFFFFFF1;
    // rom_array[39342] = 32'hFFFFFFF1;
    // rom_array[39343] = 32'hFFFFFFF1;
    // rom_array[39344] = 32'hFFFFFFF1;
    // rom_array[39345] = 32'hFFFFFFF0;
    // rom_array[39346] = 32'hFFFFFFF0;
    // rom_array[39347] = 32'hFFFFFFF0;
    // rom_array[39348] = 32'hFFFFFFF0;
    // rom_array[39349] = 32'hFFFFFFF1;
    // rom_array[39350] = 32'hFFFFFFF1;
    // rom_array[39351] = 32'hFFFFFFF1;
    // rom_array[39352] = 32'hFFFFFFF1;
    // rom_array[39353] = 32'hFFFFFFF0;
    // rom_array[39354] = 32'hFFFFFFF0;
    // rom_array[39355] = 32'hFFFFFFF0;
    // rom_array[39356] = 32'hFFFFFFF0;
    // rom_array[39357] = 32'hFFFFFFF1;
    // rom_array[39358] = 32'hFFFFFFF1;
    // rom_array[39359] = 32'hFFFFFFF1;
    // rom_array[39360] = 32'hFFFFFFF1;
    // rom_array[39361] = 32'hFFFFFFF0;
    // rom_array[39362] = 32'hFFFFFFF0;
    // rom_array[39363] = 32'hFFFFFFF0;
    // rom_array[39364] = 32'hFFFFFFF0;
    // rom_array[39365] = 32'hFFFFFFF1;
    // rom_array[39366] = 32'hFFFFFFF1;
    // rom_array[39367] = 32'hFFFFFFF1;
    // rom_array[39368] = 32'hFFFFFFF1;
    // rom_array[39369] = 32'hFFFFFFF0;
    // rom_array[39370] = 32'hFFFFFFF0;
    // rom_array[39371] = 32'hFFFFFFF0;
    // rom_array[39372] = 32'hFFFFFFF0;
    // rom_array[39373] = 32'hFFFFFFF1;
    // rom_array[39374] = 32'hFFFFFFF1;
    // rom_array[39375] = 32'hFFFFFFF1;
    // rom_array[39376] = 32'hFFFFFFF1;
    // rom_array[39377] = 32'hFFFFFFF0;
    // rom_array[39378] = 32'hFFFFFFF0;
    // rom_array[39379] = 32'hFFFFFFF0;
    // rom_array[39380] = 32'hFFFFFFF0;
    // rom_array[39381] = 32'hFFFFFFF1;
    // rom_array[39382] = 32'hFFFFFFF1;
    // rom_array[39383] = 32'hFFFFFFF1;
    // rom_array[39384] = 32'hFFFFFFF1;
    // rom_array[39385] = 32'hFFFFFFF0;
    // rom_array[39386] = 32'hFFFFFFF0;
    // rom_array[39387] = 32'hFFFFFFF0;
    // rom_array[39388] = 32'hFFFFFFF0;
    // rom_array[39389] = 32'hFFFFFFF1;
    // rom_array[39390] = 32'hFFFFFFF1;
    // rom_array[39391] = 32'hFFFFFFF1;
    // rom_array[39392] = 32'hFFFFFFF1;
    // rom_array[39393] = 32'hFFFFFFF0;
    // rom_array[39394] = 32'hFFFFFFF0;
    // rom_array[39395] = 32'hFFFFFFF0;
    // rom_array[39396] = 32'hFFFFFFF0;
    // rom_array[39397] = 32'hFFFFFFF1;
    // rom_array[39398] = 32'hFFFFFFF1;
    // rom_array[39399] = 32'hFFFFFFF1;
    // rom_array[39400] = 32'hFFFFFFF1;
    // rom_array[39401] = 32'hFFFFFFF0;
    // rom_array[39402] = 32'hFFFFFFF0;
    // rom_array[39403] = 32'hFFFFFFF0;
    // rom_array[39404] = 32'hFFFFFFF0;
    // rom_array[39405] = 32'hFFFFFFF1;
    // rom_array[39406] = 32'hFFFFFFF1;
    // rom_array[39407] = 32'hFFFFFFF1;
    // rom_array[39408] = 32'hFFFFFFF1;
    // rom_array[39409] = 32'hFFFFFFF0;
    // rom_array[39410] = 32'hFFFFFFF0;
    // rom_array[39411] = 32'hFFFFFFF0;
    // rom_array[39412] = 32'hFFFFFFF0;
    // rom_array[39413] = 32'hFFFFFFF1;
    // rom_array[39414] = 32'hFFFFFFF1;
    // rom_array[39415] = 32'hFFFFFFF1;
    // rom_array[39416] = 32'hFFFFFFF1;
    // rom_array[39417] = 32'hFFFFFFF0;
    // rom_array[39418] = 32'hFFFFFFF0;
    // rom_array[39419] = 32'hFFFFFFF0;
    // rom_array[39420] = 32'hFFFFFFF0;
    // rom_array[39421] = 32'hFFFFFFF1;
    // rom_array[39422] = 32'hFFFFFFF1;
    // rom_array[39423] = 32'hFFFFFFF1;
    // rom_array[39424] = 32'hFFFFFFF1;
    // rom_array[39425] = 32'hFFFFFFF0;
    // rom_array[39426] = 32'hFFFFFFF0;
    // rom_array[39427] = 32'hFFFFFFF0;
    // rom_array[39428] = 32'hFFFFFFF0;
    // rom_array[39429] = 32'hFFFFFFF1;
    // rom_array[39430] = 32'hFFFFFFF1;
    // rom_array[39431] = 32'hFFFFFFF1;
    // rom_array[39432] = 32'hFFFFFFF1;
    // rom_array[39433] = 32'hFFFFFFF0;
    // rom_array[39434] = 32'hFFFFFFF0;
    // rom_array[39435] = 32'hFFFFFFF0;
    // rom_array[39436] = 32'hFFFFFFF0;
    // rom_array[39437] = 32'hFFFFFFF1;
    // rom_array[39438] = 32'hFFFFFFF1;
    // rom_array[39439] = 32'hFFFFFFF1;
    // rom_array[39440] = 32'hFFFFFFF1;
    // rom_array[39441] = 32'hFFFFFFF0;
    // rom_array[39442] = 32'hFFFFFFF0;
    // rom_array[39443] = 32'hFFFFFFF0;
    // rom_array[39444] = 32'hFFFFFFF0;
    // rom_array[39445] = 32'hFFFFFFF1;
    // rom_array[39446] = 32'hFFFFFFF1;
    // rom_array[39447] = 32'hFFFFFFF1;
    // rom_array[39448] = 32'hFFFFFFF1;
    // rom_array[39449] = 32'hFFFFFFF0;
    // rom_array[39450] = 32'hFFFFFFF0;
    // rom_array[39451] = 32'hFFFFFFF0;
    // rom_array[39452] = 32'hFFFFFFF0;
    // rom_array[39453] = 32'hFFFFFFF1;
    // rom_array[39454] = 32'hFFFFFFF1;
    // rom_array[39455] = 32'hFFFFFFF1;
    // rom_array[39456] = 32'hFFFFFFF1;
    // rom_array[39457] = 32'hFFFFFFF0;
    // rom_array[39458] = 32'hFFFFFFF0;
    // rom_array[39459] = 32'hFFFFFFF0;
    // rom_array[39460] = 32'hFFFFFFF0;
    // rom_array[39461] = 32'hFFFFFFF1;
    // rom_array[39462] = 32'hFFFFFFF1;
    // rom_array[39463] = 32'hFFFFFFF1;
    // rom_array[39464] = 32'hFFFFFFF1;
    // rom_array[39465] = 32'hFFFFFFF1;
    // rom_array[39466] = 32'hFFFFFFF1;
    // rom_array[39467] = 32'hFFFFFFF1;
    // rom_array[39468] = 32'hFFFFFFF1;
    // rom_array[39469] = 32'hFFFFFFF1;
    // rom_array[39470] = 32'hFFFFFFF1;
    // rom_array[39471] = 32'hFFFFFFF1;
    // rom_array[39472] = 32'hFFFFFFF1;
    // rom_array[39473] = 32'hFFFFFFF1;
    // rom_array[39474] = 32'hFFFFFFF1;
    // rom_array[39475] = 32'hFFFFFFF1;
    // rom_array[39476] = 32'hFFFFFFF1;
    // rom_array[39477] = 32'hFFFFFFF1;
    // rom_array[39478] = 32'hFFFFFFF1;
    // rom_array[39479] = 32'hFFFFFFF1;
    // rom_array[39480] = 32'hFFFFFFF1;
    // rom_array[39481] = 32'hFFFFFFF1;
    // rom_array[39482] = 32'hFFFFFFF1;
    // rom_array[39483] = 32'hFFFFFFF1;
    // rom_array[39484] = 32'hFFFFFFF1;
    // rom_array[39485] = 32'hFFFFFFF0;
    // rom_array[39486] = 32'hFFFFFFF0;
    // rom_array[39487] = 32'hFFFFFFF0;
    // rom_array[39488] = 32'hFFFFFFF0;
    // rom_array[39489] = 32'hFFFFFFF1;
    // rom_array[39490] = 32'hFFFFFFF1;
    // rom_array[39491] = 32'hFFFFFFF1;
    // rom_array[39492] = 32'hFFFFFFF1;
    // rom_array[39493] = 32'hFFFFFFF0;
    // rom_array[39494] = 32'hFFFFFFF0;
    // rom_array[39495] = 32'hFFFFFFF0;
    // rom_array[39496] = 32'hFFFFFFF0;
    // rom_array[39497] = 32'hFFFFFFF1;
    // rom_array[39498] = 32'hFFFFFFF1;
    // rom_array[39499] = 32'hFFFFFFF1;
    // rom_array[39500] = 32'hFFFFFFF1;
    // rom_array[39501] = 32'hFFFFFFF1;
    // rom_array[39502] = 32'hFFFFFFF1;
    // rom_array[39503] = 32'hFFFFFFF1;
    // rom_array[39504] = 32'hFFFFFFF1;
    // rom_array[39505] = 32'hFFFFFFF1;
    // rom_array[39506] = 32'hFFFFFFF1;
    // rom_array[39507] = 32'hFFFFFFF1;
    // rom_array[39508] = 32'hFFFFFFF1;
    // rom_array[39509] = 32'hFFFFFFF1;
    // rom_array[39510] = 32'hFFFFFFF1;
    // rom_array[39511] = 32'hFFFFFFF1;
    // rom_array[39512] = 32'hFFFFFFF1;
    // rom_array[39513] = 32'hFFFFFFF1;
    // rom_array[39514] = 32'hFFFFFFF1;
    // rom_array[39515] = 32'hFFFFFFF1;
    // rom_array[39516] = 32'hFFFFFFF1;
    // rom_array[39517] = 32'hFFFFFFF0;
    // rom_array[39518] = 32'hFFFFFFF0;
    // rom_array[39519] = 32'hFFFFFFF0;
    // rom_array[39520] = 32'hFFFFFFF0;
    // rom_array[39521] = 32'hFFFFFFF1;
    // rom_array[39522] = 32'hFFFFFFF1;
    // rom_array[39523] = 32'hFFFFFFF1;
    // rom_array[39524] = 32'hFFFFFFF1;
    // rom_array[39525] = 32'hFFFFFFF0;
    // rom_array[39526] = 32'hFFFFFFF0;
    // rom_array[39527] = 32'hFFFFFFF0;
    // rom_array[39528] = 32'hFFFFFFF0;
    // rom_array[39529] = 32'hFFFFFFF1;
    // rom_array[39530] = 32'hFFFFFFF1;
    // rom_array[39531] = 32'hFFFFFFF1;
    // rom_array[39532] = 32'hFFFFFFF1;
    // rom_array[39533] = 32'hFFFFFFF0;
    // rom_array[39534] = 32'hFFFFFFF0;
    // rom_array[39535] = 32'hFFFFFFF0;
    // rom_array[39536] = 32'hFFFFFFF0;
    // rom_array[39537] = 32'hFFFFFFF1;
    // rom_array[39538] = 32'hFFFFFFF1;
    // rom_array[39539] = 32'hFFFFFFF1;
    // rom_array[39540] = 32'hFFFFFFF1;
    // rom_array[39541] = 32'hFFFFFFF0;
    // rom_array[39542] = 32'hFFFFFFF0;
    // rom_array[39543] = 32'hFFFFFFF0;
    // rom_array[39544] = 32'hFFFFFFF0;
    // rom_array[39545] = 32'hFFFFFFF1;
    // rom_array[39546] = 32'hFFFFFFF1;
    // rom_array[39547] = 32'hFFFFFFF1;
    // rom_array[39548] = 32'hFFFFFFF1;
    // rom_array[39549] = 32'hFFFFFFF0;
    // rom_array[39550] = 32'hFFFFFFF0;
    // rom_array[39551] = 32'hFFFFFFF0;
    // rom_array[39552] = 32'hFFFFFFF0;
    // rom_array[39553] = 32'hFFFFFFF1;
    // rom_array[39554] = 32'hFFFFFFF1;
    // rom_array[39555] = 32'hFFFFFFF1;
    // rom_array[39556] = 32'hFFFFFFF1;
    // rom_array[39557] = 32'hFFFFFFF0;
    // rom_array[39558] = 32'hFFFFFFF0;
    // rom_array[39559] = 32'hFFFFFFF0;
    // rom_array[39560] = 32'hFFFFFFF0;
    // rom_array[39561] = 32'hFFFFFFF1;
    // rom_array[39562] = 32'hFFFFFFF1;
    // rom_array[39563] = 32'hFFFFFFF1;
    // rom_array[39564] = 32'hFFFFFFF1;
    // rom_array[39565] = 32'hFFFFFFF0;
    // rom_array[39566] = 32'hFFFFFFF0;
    // rom_array[39567] = 32'hFFFFFFF0;
    // rom_array[39568] = 32'hFFFFFFF0;
    // rom_array[39569] = 32'hFFFFFFF1;
    // rom_array[39570] = 32'hFFFFFFF1;
    // rom_array[39571] = 32'hFFFFFFF1;
    // rom_array[39572] = 32'hFFFFFFF1;
    // rom_array[39573] = 32'hFFFFFFF0;
    // rom_array[39574] = 32'hFFFFFFF0;
    // rom_array[39575] = 32'hFFFFFFF0;
    // rom_array[39576] = 32'hFFFFFFF0;
    // rom_array[39577] = 32'hFFFFFFF1;
    // rom_array[39578] = 32'hFFFFFFF1;
    // rom_array[39579] = 32'hFFFFFFF1;
    // rom_array[39580] = 32'hFFFFFFF1;
    // rom_array[39581] = 32'hFFFFFFF0;
    // rom_array[39582] = 32'hFFFFFFF0;
    // rom_array[39583] = 32'hFFFFFFF1;
    // rom_array[39584] = 32'hFFFFFFF1;
    // rom_array[39585] = 32'hFFFFFFF1;
    // rom_array[39586] = 32'hFFFFFFF1;
    // rom_array[39587] = 32'hFFFFFFF1;
    // rom_array[39588] = 32'hFFFFFFF1;
    // rom_array[39589] = 32'hFFFFFFF0;
    // rom_array[39590] = 32'hFFFFFFF0;
    // rom_array[39591] = 32'hFFFFFFF1;
    // rom_array[39592] = 32'hFFFFFFF1;
    // rom_array[39593] = 32'hFFFFFFF1;
    // rom_array[39594] = 32'hFFFFFFF1;
    // rom_array[39595] = 32'hFFFFFFF1;
    // rom_array[39596] = 32'hFFFFFFF1;
    // rom_array[39597] = 32'hFFFFFFF1;
    // rom_array[39598] = 32'hFFFFFFF1;
    // rom_array[39599] = 32'hFFFFFFF1;
    // rom_array[39600] = 32'hFFFFFFF1;
    // rom_array[39601] = 32'hFFFFFFF1;
    // rom_array[39602] = 32'hFFFFFFF1;
    // rom_array[39603] = 32'hFFFFFFF1;
    // rom_array[39604] = 32'hFFFFFFF1;
    // rom_array[39605] = 32'hFFFFFFF1;
    // rom_array[39606] = 32'hFFFFFFF1;
    // rom_array[39607] = 32'hFFFFFFF1;
    // rom_array[39608] = 32'hFFFFFFF1;
    // rom_array[39609] = 32'hFFFFFFF0;
    // rom_array[39610] = 32'hFFFFFFF0;
    // rom_array[39611] = 32'hFFFFFFF1;
    // rom_array[39612] = 32'hFFFFFFF1;
    // rom_array[39613] = 32'hFFFFFFF0;
    // rom_array[39614] = 32'hFFFFFFF0;
    // rom_array[39615] = 32'hFFFFFFF1;
    // rom_array[39616] = 32'hFFFFFFF1;
    // rom_array[39617] = 32'hFFFFFFF0;
    // rom_array[39618] = 32'hFFFFFFF0;
    // rom_array[39619] = 32'hFFFFFFF1;
    // rom_array[39620] = 32'hFFFFFFF1;
    // rom_array[39621] = 32'hFFFFFFF0;
    // rom_array[39622] = 32'hFFFFFFF0;
    // rom_array[39623] = 32'hFFFFFFF1;
    // rom_array[39624] = 32'hFFFFFFF1;
    // rom_array[39625] = 32'hFFFFFFF0;
    // rom_array[39626] = 32'hFFFFFFF0;
    // rom_array[39627] = 32'hFFFFFFF0;
    // rom_array[39628] = 32'hFFFFFFF0;
    // rom_array[39629] = 32'hFFFFFFF1;
    // rom_array[39630] = 32'hFFFFFFF1;
    // rom_array[39631] = 32'hFFFFFFF1;
    // rom_array[39632] = 32'hFFFFFFF1;
    // rom_array[39633] = 32'hFFFFFFF0;
    // rom_array[39634] = 32'hFFFFFFF0;
    // rom_array[39635] = 32'hFFFFFFF0;
    // rom_array[39636] = 32'hFFFFFFF0;
    // rom_array[39637] = 32'hFFFFFFF1;
    // rom_array[39638] = 32'hFFFFFFF1;
    // rom_array[39639] = 32'hFFFFFFF1;
    // rom_array[39640] = 32'hFFFFFFF1;
    // rom_array[39641] = 32'hFFFFFFF0;
    // rom_array[39642] = 32'hFFFFFFF0;
    // rom_array[39643] = 32'hFFFFFFF0;
    // rom_array[39644] = 32'hFFFFFFF0;
    // rom_array[39645] = 32'hFFFFFFF1;
    // rom_array[39646] = 32'hFFFFFFF1;
    // rom_array[39647] = 32'hFFFFFFF1;
    // rom_array[39648] = 32'hFFFFFFF1;
    // rom_array[39649] = 32'hFFFFFFF0;
    // rom_array[39650] = 32'hFFFFFFF0;
    // rom_array[39651] = 32'hFFFFFFF0;
    // rom_array[39652] = 32'hFFFFFFF0;
    // rom_array[39653] = 32'hFFFFFFF1;
    // rom_array[39654] = 32'hFFFFFFF1;
    // rom_array[39655] = 32'hFFFFFFF1;
    // rom_array[39656] = 32'hFFFFFFF1;
    // rom_array[39657] = 32'hFFFFFFF0;
    // rom_array[39658] = 32'hFFFFFFF0;
    // rom_array[39659] = 32'hFFFFFFF0;
    // rom_array[39660] = 32'hFFFFFFF0;
    // rom_array[39661] = 32'hFFFFFFF1;
    // rom_array[39662] = 32'hFFFFFFF1;
    // rom_array[39663] = 32'hFFFFFFF1;
    // rom_array[39664] = 32'hFFFFFFF1;
    // rom_array[39665] = 32'hFFFFFFF0;
    // rom_array[39666] = 32'hFFFFFFF0;
    // rom_array[39667] = 32'hFFFFFFF0;
    // rom_array[39668] = 32'hFFFFFFF0;
    // rom_array[39669] = 32'hFFFFFFF1;
    // rom_array[39670] = 32'hFFFFFFF1;
    // rom_array[39671] = 32'hFFFFFFF1;
    // rom_array[39672] = 32'hFFFFFFF1;
    // rom_array[39673] = 32'hFFFFFFF1;
    // rom_array[39674] = 32'hFFFFFFF1;
    // rom_array[39675] = 32'hFFFFFFF1;
    // rom_array[39676] = 32'hFFFFFFF1;
    // rom_array[39677] = 32'hFFFFFFF1;
    // rom_array[39678] = 32'hFFFFFFF1;
    // rom_array[39679] = 32'hFFFFFFF1;
    // rom_array[39680] = 32'hFFFFFFF1;
    // rom_array[39681] = 32'hFFFFFFF1;
    // rom_array[39682] = 32'hFFFFFFF1;
    // rom_array[39683] = 32'hFFFFFFF1;
    // rom_array[39684] = 32'hFFFFFFF1;
    // rom_array[39685] = 32'hFFFFFFF1;
    // rom_array[39686] = 32'hFFFFFFF1;
    // rom_array[39687] = 32'hFFFFFFF1;
    // rom_array[39688] = 32'hFFFFFFF1;
    // rom_array[39689] = 32'hFFFFFFF1;
    // rom_array[39690] = 32'hFFFFFFF1;
    // rom_array[39691] = 32'hFFFFFFF1;
    // rom_array[39692] = 32'hFFFFFFF1;
    // rom_array[39693] = 32'hFFFFFFF1;
    // rom_array[39694] = 32'hFFFFFFF1;
    // rom_array[39695] = 32'hFFFFFFF1;
    // rom_array[39696] = 32'hFFFFFFF1;
    // rom_array[39697] = 32'hFFFFFFF1;
    // rom_array[39698] = 32'hFFFFFFF1;
    // rom_array[39699] = 32'hFFFFFFF1;
    // rom_array[39700] = 32'hFFFFFFF1;
    // rom_array[39701] = 32'hFFFFFFF1;
    // rom_array[39702] = 32'hFFFFFFF1;
    // rom_array[39703] = 32'hFFFFFFF1;
    // rom_array[39704] = 32'hFFFFFFF1;
    // rom_array[39705] = 32'hFFFFFFF1;
    // rom_array[39706] = 32'hFFFFFFF1;
    // rom_array[39707] = 32'hFFFFFFF1;
    // rom_array[39708] = 32'hFFFFFFF1;
    // rom_array[39709] = 32'hFFFFFFF1;
    // rom_array[39710] = 32'hFFFFFFF1;
    // rom_array[39711] = 32'hFFFFFFF1;
    // rom_array[39712] = 32'hFFFFFFF1;
    // rom_array[39713] = 32'hFFFFFFF1;
    // rom_array[39714] = 32'hFFFFFFF1;
    // rom_array[39715] = 32'hFFFFFFF1;
    // rom_array[39716] = 32'hFFFFFFF1;
    // rom_array[39717] = 32'hFFFFFFF1;
    // rom_array[39718] = 32'hFFFFFFF1;
    // rom_array[39719] = 32'hFFFFFFF1;
    // rom_array[39720] = 32'hFFFFFFF1;
    // rom_array[39721] = 32'hFFFFFFF1;
    // rom_array[39722] = 32'hFFFFFFF1;
    // rom_array[39723] = 32'hFFFFFFF1;
    // rom_array[39724] = 32'hFFFFFFF1;
    // rom_array[39725] = 32'hFFFFFFF1;
    // rom_array[39726] = 32'hFFFFFFF1;
    // rom_array[39727] = 32'hFFFFFFF1;
    // rom_array[39728] = 32'hFFFFFFF1;
    // rom_array[39729] = 32'hFFFFFFF1;
    // rom_array[39730] = 32'hFFFFFFF1;
    // rom_array[39731] = 32'hFFFFFFF1;
    // rom_array[39732] = 32'hFFFFFFF1;
    // rom_array[39733] = 32'hFFFFFFF1;
    // rom_array[39734] = 32'hFFFFFFF1;
    // rom_array[39735] = 32'hFFFFFFF1;
    // rom_array[39736] = 32'hFFFFFFF1;
    // rom_array[39737] = 32'hFFFFFFF1;
    // rom_array[39738] = 32'hFFFFFFF1;
    // rom_array[39739] = 32'hFFFFFFF1;
    // rom_array[39740] = 32'hFFFFFFF1;
    // rom_array[39741] = 32'hFFFFFFF1;
    // rom_array[39742] = 32'hFFFFFFF1;
    // rom_array[39743] = 32'hFFFFFFF1;
    // rom_array[39744] = 32'hFFFFFFF1;
    // rom_array[39745] = 32'hFFFFFFF1;
    // rom_array[39746] = 32'hFFFFFFF1;
    // rom_array[39747] = 32'hFFFFFFF1;
    // rom_array[39748] = 32'hFFFFFFF1;
    // rom_array[39749] = 32'hFFFFFFF1;
    // rom_array[39750] = 32'hFFFFFFF1;
    // rom_array[39751] = 32'hFFFFFFF1;
    // rom_array[39752] = 32'hFFFFFFF1;
    // rom_array[39753] = 32'hFFFFFFF1;
    // rom_array[39754] = 32'hFFFFFFF1;
    // rom_array[39755] = 32'hFFFFFFF1;
    // rom_array[39756] = 32'hFFFFFFF1;
    // rom_array[39757] = 32'hFFFFFFF1;
    // rom_array[39758] = 32'hFFFFFFF1;
    // rom_array[39759] = 32'hFFFFFFF1;
    // rom_array[39760] = 32'hFFFFFFF1;
    // rom_array[39761] = 32'hFFFFFFF1;
    // rom_array[39762] = 32'hFFFFFFF1;
    // rom_array[39763] = 32'hFFFFFFF1;
    // rom_array[39764] = 32'hFFFFFFF1;
    // rom_array[39765] = 32'hFFFFFFF1;
    // rom_array[39766] = 32'hFFFFFFF1;
    // rom_array[39767] = 32'hFFFFFFF1;
    // rom_array[39768] = 32'hFFFFFFF1;
    // rom_array[39769] = 32'hFFFFFFF1;
    // rom_array[39770] = 32'hFFFFFFF1;
    // rom_array[39771] = 32'hFFFFFFF1;
    // rom_array[39772] = 32'hFFFFFFF1;
    // rom_array[39773] = 32'hFFFFFFF1;
    // rom_array[39774] = 32'hFFFFFFF1;
    // rom_array[39775] = 32'hFFFFFFF1;
    // rom_array[39776] = 32'hFFFFFFF1;
    // rom_array[39777] = 32'hFFFFFFF1;
    // rom_array[39778] = 32'hFFFFFFF1;
    // rom_array[39779] = 32'hFFFFFFF1;
    // rom_array[39780] = 32'hFFFFFFF1;
    // rom_array[39781] = 32'hFFFFFFF1;
    // rom_array[39782] = 32'hFFFFFFF1;
    // rom_array[39783] = 32'hFFFFFFF1;
    // rom_array[39784] = 32'hFFFFFFF1;
    // rom_array[39785] = 32'hFFFFFFF1;
    // rom_array[39786] = 32'hFFFFFFF1;
    // rom_array[39787] = 32'hFFFFFFF1;
    // rom_array[39788] = 32'hFFFFFFF1;
    // rom_array[39789] = 32'hFFFFFFF1;
    // rom_array[39790] = 32'hFFFFFFF1;
    // rom_array[39791] = 32'hFFFFFFF1;
    // rom_array[39792] = 32'hFFFFFFF1;
    // rom_array[39793] = 32'hFFFFFFF1;
    // rom_array[39794] = 32'hFFFFFFF1;
    // rom_array[39795] = 32'hFFFFFFF1;
    // rom_array[39796] = 32'hFFFFFFF1;
    // rom_array[39797] = 32'hFFFFFFF1;
    // rom_array[39798] = 32'hFFFFFFF1;
    // rom_array[39799] = 32'hFFFFFFF1;
    // rom_array[39800] = 32'hFFFFFFF1;
    // rom_array[39801] = 32'hFFFFFFF1;
    // rom_array[39802] = 32'hFFFFFFF1;
    // rom_array[39803] = 32'hFFFFFFF1;
    // rom_array[39804] = 32'hFFFFFFF1;
    // rom_array[39805] = 32'hFFFFFFF1;
    // rom_array[39806] = 32'hFFFFFFF1;
    // rom_array[39807] = 32'hFFFFFFF1;
    // rom_array[39808] = 32'hFFFFFFF1;
    // rom_array[39809] = 32'hFFFFFFF1;
    // rom_array[39810] = 32'hFFFFFFF1;
    // rom_array[39811] = 32'hFFFFFFF1;
    // rom_array[39812] = 32'hFFFFFFF1;
    // rom_array[39813] = 32'hFFFFFFF1;
    // rom_array[39814] = 32'hFFFFFFF1;
    // rom_array[39815] = 32'hFFFFFFF1;
    // rom_array[39816] = 32'hFFFFFFF1;
    // rom_array[39817] = 32'hFFFFFFF1;
    // rom_array[39818] = 32'hFFFFFFF1;
    // rom_array[39819] = 32'hFFFFFFF1;
    // rom_array[39820] = 32'hFFFFFFF1;
    // rom_array[39821] = 32'hFFFFFFF1;
    // rom_array[39822] = 32'hFFFFFFF1;
    // rom_array[39823] = 32'hFFFFFFF1;
    // rom_array[39824] = 32'hFFFFFFF1;
    // rom_array[39825] = 32'hFFFFFFF1;
    // rom_array[39826] = 32'hFFFFFFF1;
    // rom_array[39827] = 32'hFFFFFFF1;
    // rom_array[39828] = 32'hFFFFFFF1;
    // rom_array[39829] = 32'hFFFFFFF1;
    // rom_array[39830] = 32'hFFFFFFF1;
    // rom_array[39831] = 32'hFFFFFFF1;
    // rom_array[39832] = 32'hFFFFFFF1;
    // rom_array[39833] = 32'hFFFFFFF1;
    // rom_array[39834] = 32'hFFFFFFF1;
    // rom_array[39835] = 32'hFFFFFFF1;
    // rom_array[39836] = 32'hFFFFFFF1;
    // rom_array[39837] = 32'hFFFFFFF1;
    // rom_array[39838] = 32'hFFFFFFF1;
    // rom_array[39839] = 32'hFFFFFFF1;
    // rom_array[39840] = 32'hFFFFFFF1;
    // rom_array[39841] = 32'hFFFFFFF1;
    // rom_array[39842] = 32'hFFFFFFF1;
    // rom_array[39843] = 32'hFFFFFFF1;
    // rom_array[39844] = 32'hFFFFFFF1;
    // rom_array[39845] = 32'hFFFFFFF1;
    // rom_array[39846] = 32'hFFFFFFF1;
    // rom_array[39847] = 32'hFFFFFFF1;
    // rom_array[39848] = 32'hFFFFFFF1;
    // rom_array[39849] = 32'hFFFFFFF0;
    // rom_array[39850] = 32'hFFFFFFF0;
    // rom_array[39851] = 32'hFFFFFFF1;
    // rom_array[39852] = 32'hFFFFFFF1;
    // rom_array[39853] = 32'hFFFFFFF0;
    // rom_array[39854] = 32'hFFFFFFF0;
    // rom_array[39855] = 32'hFFFFFFF1;
    // rom_array[39856] = 32'hFFFFFFF1;
    // rom_array[39857] = 32'hFFFFFFF0;
    // rom_array[39858] = 32'hFFFFFFF0;
    // rom_array[39859] = 32'hFFFFFFF1;
    // rom_array[39860] = 32'hFFFFFFF1;
    // rom_array[39861] = 32'hFFFFFFF0;
    // rom_array[39862] = 32'hFFFFFFF0;
    // rom_array[39863] = 32'hFFFFFFF1;
    // rom_array[39864] = 32'hFFFFFFF1;
    // rom_array[39865] = 32'hFFFFFFF0;
    // rom_array[39866] = 32'hFFFFFFF0;
    // rom_array[39867] = 32'hFFFFFFF1;
    // rom_array[39868] = 32'hFFFFFFF1;
    // rom_array[39869] = 32'hFFFFFFF0;
    // rom_array[39870] = 32'hFFFFFFF0;
    // rom_array[39871] = 32'hFFFFFFF1;
    // rom_array[39872] = 32'hFFFFFFF1;
    // rom_array[39873] = 32'hFFFFFFF0;
    // rom_array[39874] = 32'hFFFFFFF0;
    // rom_array[39875] = 32'hFFFFFFF1;
    // rom_array[39876] = 32'hFFFFFFF1;
    // rom_array[39877] = 32'hFFFFFFF0;
    // rom_array[39878] = 32'hFFFFFFF0;
    // rom_array[39879] = 32'hFFFFFFF1;
    // rom_array[39880] = 32'hFFFFFFF1;
    // rom_array[39881] = 32'hFFFFFFF0;
    // rom_array[39882] = 32'hFFFFFFF0;
    // rom_array[39883] = 32'hFFFFFFF1;
    // rom_array[39884] = 32'hFFFFFFF1;
    // rom_array[39885] = 32'hFFFFFFF0;
    // rom_array[39886] = 32'hFFFFFFF0;
    // rom_array[39887] = 32'hFFFFFFF1;
    // rom_array[39888] = 32'hFFFFFFF1;
    // rom_array[39889] = 32'hFFFFFFF0;
    // rom_array[39890] = 32'hFFFFFFF0;
    // rom_array[39891] = 32'hFFFFFFF1;
    // rom_array[39892] = 32'hFFFFFFF1;
    // rom_array[39893] = 32'hFFFFFFF0;
    // rom_array[39894] = 32'hFFFFFFF0;
    // rom_array[39895] = 32'hFFFFFFF1;
    // rom_array[39896] = 32'hFFFFFFF1;
    // rom_array[39897] = 32'hFFFFFFF0;
    // rom_array[39898] = 32'hFFFFFFF0;
    // rom_array[39899] = 32'hFFFFFFF1;
    // rom_array[39900] = 32'hFFFFFFF1;
    // rom_array[39901] = 32'hFFFFFFF0;
    // rom_array[39902] = 32'hFFFFFFF0;
    // rom_array[39903] = 32'hFFFFFFF1;
    // rom_array[39904] = 32'hFFFFFFF1;
    // rom_array[39905] = 32'hFFFFFFF0;
    // rom_array[39906] = 32'hFFFFFFF0;
    // rom_array[39907] = 32'hFFFFFFF1;
    // rom_array[39908] = 32'hFFFFFFF1;
    // rom_array[39909] = 32'hFFFFFFF0;
    // rom_array[39910] = 32'hFFFFFFF0;
    // rom_array[39911] = 32'hFFFFFFF1;
    // rom_array[39912] = 32'hFFFFFFF1;
    // rom_array[39913] = 32'hFFFFFFF1;
    // rom_array[39914] = 32'hFFFFFFF1;
    // rom_array[39915] = 32'hFFFFFFF1;
    // rom_array[39916] = 32'hFFFFFFF1;
    // rom_array[39917] = 32'hFFFFFFF1;
    // rom_array[39918] = 32'hFFFFFFF1;
    // rom_array[39919] = 32'hFFFFFFF1;
    // rom_array[39920] = 32'hFFFFFFF1;
    // rom_array[39921] = 32'hFFFFFFF1;
    // rom_array[39922] = 32'hFFFFFFF1;
    // rom_array[39923] = 32'hFFFFFFF1;
    // rom_array[39924] = 32'hFFFFFFF1;
    // rom_array[39925] = 32'hFFFFFFF1;
    // rom_array[39926] = 32'hFFFFFFF1;
    // rom_array[39927] = 32'hFFFFFFF1;
    // rom_array[39928] = 32'hFFFFFFF1;
    // rom_array[39929] = 32'hFFFFFFF1;
    // rom_array[39930] = 32'hFFFFFFF1;
    // rom_array[39931] = 32'hFFFFFFF1;
    // rom_array[39932] = 32'hFFFFFFF1;
    // rom_array[39933] = 32'hFFFFFFF1;
    // rom_array[39934] = 32'hFFFFFFF1;
    // rom_array[39935] = 32'hFFFFFFF1;
    // rom_array[39936] = 32'hFFFFFFF1;
    // rom_array[39937] = 32'hFFFFFFF1;
    // rom_array[39938] = 32'hFFFFFFF1;
    // rom_array[39939] = 32'hFFFFFFF1;
    // rom_array[39940] = 32'hFFFFFFF1;
    // rom_array[39941] = 32'hFFFFFFF1;
    // rom_array[39942] = 32'hFFFFFFF1;
    // rom_array[39943] = 32'hFFFFFFF1;
    // rom_array[39944] = 32'hFFFFFFF1;
    // rom_array[39945] = 32'hFFFFFFF0;
    // rom_array[39946] = 32'hFFFFFFF0;
    // rom_array[39947] = 32'hFFFFFFF0;
    // rom_array[39948] = 32'hFFFFFFF0;
    // rom_array[39949] = 32'hFFFFFFF1;
    // rom_array[39950] = 32'hFFFFFFF1;
    // rom_array[39951] = 32'hFFFFFFF1;
    // rom_array[39952] = 32'hFFFFFFF1;
    // rom_array[39953] = 32'hFFFFFFF0;
    // rom_array[39954] = 32'hFFFFFFF0;
    // rom_array[39955] = 32'hFFFFFFF0;
    // rom_array[39956] = 32'hFFFFFFF0;
    // rom_array[39957] = 32'hFFFFFFF1;
    // rom_array[39958] = 32'hFFFFFFF1;
    // rom_array[39959] = 32'hFFFFFFF1;
    // rom_array[39960] = 32'hFFFFFFF1;
    // rom_array[39961] = 32'hFFFFFFF0;
    // rom_array[39962] = 32'hFFFFFFF0;
    // rom_array[39963] = 32'hFFFFFFF0;
    // rom_array[39964] = 32'hFFFFFFF0;
    // rom_array[39965] = 32'hFFFFFFF1;
    // rom_array[39966] = 32'hFFFFFFF1;
    // rom_array[39967] = 32'hFFFFFFF1;
    // rom_array[39968] = 32'hFFFFFFF1;
    // rom_array[39969] = 32'hFFFFFFF0;
    // rom_array[39970] = 32'hFFFFFFF0;
    // rom_array[39971] = 32'hFFFFFFF0;
    // rom_array[39972] = 32'hFFFFFFF0;
    // rom_array[39973] = 32'hFFFFFFF1;
    // rom_array[39974] = 32'hFFFFFFF1;
    // rom_array[39975] = 32'hFFFFFFF1;
    // rom_array[39976] = 32'hFFFFFFF1;
    // rom_array[39977] = 32'hFFFFFFF0;
    // rom_array[39978] = 32'hFFFFFFF0;
    // rom_array[39979] = 32'hFFFFFFF0;
    // rom_array[39980] = 32'hFFFFFFF0;
    // rom_array[39981] = 32'hFFFFFFF1;
    // rom_array[39982] = 32'hFFFFFFF1;
    // rom_array[39983] = 32'hFFFFFFF1;
    // rom_array[39984] = 32'hFFFFFFF1;
    // rom_array[39985] = 32'hFFFFFFF0;
    // rom_array[39986] = 32'hFFFFFFF0;
    // rom_array[39987] = 32'hFFFFFFF0;
    // rom_array[39988] = 32'hFFFFFFF0;
    // rom_array[39989] = 32'hFFFFFFF1;
    // rom_array[39990] = 32'hFFFFFFF1;
    // rom_array[39991] = 32'hFFFFFFF1;
    // rom_array[39992] = 32'hFFFFFFF1;
    // rom_array[39993] = 32'hFFFFFFF1;
    // rom_array[39994] = 32'hFFFFFFF1;
    // rom_array[39995] = 32'hFFFFFFF1;
    // rom_array[39996] = 32'hFFFFFFF1;
    // rom_array[39997] = 32'hFFFFFFF0;
    // rom_array[39998] = 32'hFFFFFFF0;
    // rom_array[39999] = 32'hFFFFFFF0;
    // rom_array[40000] = 32'hFFFFFFF0;
    // rom_array[40001] = 32'hFFFFFFF1;
    // rom_array[40002] = 32'hFFFFFFF1;
    // rom_array[40003] = 32'hFFFFFFF1;
    // rom_array[40004] = 32'hFFFFFFF1;
    // rom_array[40005] = 32'hFFFFFFF0;
    // rom_array[40006] = 32'hFFFFFFF0;
    // rom_array[40007] = 32'hFFFFFFF0;
    // rom_array[40008] = 32'hFFFFFFF0;
    // rom_array[40009] = 32'hFFFFFFF0;
    // rom_array[40010] = 32'hFFFFFFF0;
    // rom_array[40011] = 32'hFFFFFFF0;
    // rom_array[40012] = 32'hFFFFFFF0;
    // rom_array[40013] = 32'hFFFFFFF1;
    // rom_array[40014] = 32'hFFFFFFF1;
    // rom_array[40015] = 32'hFFFFFFF1;
    // rom_array[40016] = 32'hFFFFFFF1;
    // rom_array[40017] = 32'hFFFFFFF0;
    // rom_array[40018] = 32'hFFFFFFF0;
    // rom_array[40019] = 32'hFFFFFFF0;
    // rom_array[40020] = 32'hFFFFFFF0;
    // rom_array[40021] = 32'hFFFFFFF1;
    // rom_array[40022] = 32'hFFFFFFF1;
    // rom_array[40023] = 32'hFFFFFFF1;
    // rom_array[40024] = 32'hFFFFFFF1;
    // rom_array[40025] = 32'hFFFFFFF0;
    // rom_array[40026] = 32'hFFFFFFF0;
    // rom_array[40027] = 32'hFFFFFFF0;
    // rom_array[40028] = 32'hFFFFFFF0;
    // rom_array[40029] = 32'hFFFFFFF1;
    // rom_array[40030] = 32'hFFFFFFF1;
    // rom_array[40031] = 32'hFFFFFFF1;
    // rom_array[40032] = 32'hFFFFFFF1;
    // rom_array[40033] = 32'hFFFFFFF0;
    // rom_array[40034] = 32'hFFFFFFF0;
    // rom_array[40035] = 32'hFFFFFFF0;
    // rom_array[40036] = 32'hFFFFFFF0;
    // rom_array[40037] = 32'hFFFFFFF1;
    // rom_array[40038] = 32'hFFFFFFF1;
    // rom_array[40039] = 32'hFFFFFFF1;
    // rom_array[40040] = 32'hFFFFFFF1;
    // rom_array[40041] = 32'hFFFFFFF0;
    // rom_array[40042] = 32'hFFFFFFF0;
    // rom_array[40043] = 32'hFFFFFFF1;
    // rom_array[40044] = 32'hFFFFFFF1;
    // rom_array[40045] = 32'hFFFFFFF0;
    // rom_array[40046] = 32'hFFFFFFF0;
    // rom_array[40047] = 32'hFFFFFFF1;
    // rom_array[40048] = 32'hFFFFFFF1;
    // rom_array[40049] = 32'hFFFFFFF0;
    // rom_array[40050] = 32'hFFFFFFF0;
    // rom_array[40051] = 32'hFFFFFFF1;
    // rom_array[40052] = 32'hFFFFFFF1;
    // rom_array[40053] = 32'hFFFFFFF0;
    // rom_array[40054] = 32'hFFFFFFF0;
    // rom_array[40055] = 32'hFFFFFFF1;
    // rom_array[40056] = 32'hFFFFFFF1;
    // rom_array[40057] = 32'hFFFFFFF0;
    // rom_array[40058] = 32'hFFFFFFF0;
    // rom_array[40059] = 32'hFFFFFFF1;
    // rom_array[40060] = 32'hFFFFFFF1;
    // rom_array[40061] = 32'hFFFFFFF1;
    // rom_array[40062] = 32'hFFFFFFF1;
    // rom_array[40063] = 32'hFFFFFFF1;
    // rom_array[40064] = 32'hFFFFFFF1;
    // rom_array[40065] = 32'hFFFFFFF0;
    // rom_array[40066] = 32'hFFFFFFF0;
    // rom_array[40067] = 32'hFFFFFFF1;
    // rom_array[40068] = 32'hFFFFFFF1;
    // rom_array[40069] = 32'hFFFFFFF1;
    // rom_array[40070] = 32'hFFFFFFF1;
    // rom_array[40071] = 32'hFFFFFFF1;
    // rom_array[40072] = 32'hFFFFFFF1;
    // rom_array[40073] = 32'hFFFFFFF0;
    // rom_array[40074] = 32'hFFFFFFF0;
    // rom_array[40075] = 32'hFFFFFFF0;
    // rom_array[40076] = 32'hFFFFFFF0;
    // rom_array[40077] = 32'hFFFFFFF1;
    // rom_array[40078] = 32'hFFFFFFF1;
    // rom_array[40079] = 32'hFFFFFFF1;
    // rom_array[40080] = 32'hFFFFFFF1;
    // rom_array[40081] = 32'hFFFFFFF0;
    // rom_array[40082] = 32'hFFFFFFF0;
    // rom_array[40083] = 32'hFFFFFFF0;
    // rom_array[40084] = 32'hFFFFFFF0;
    // rom_array[40085] = 32'hFFFFFFF1;
    // rom_array[40086] = 32'hFFFFFFF1;
    // rom_array[40087] = 32'hFFFFFFF1;
    // rom_array[40088] = 32'hFFFFFFF1;
    // rom_array[40089] = 32'hFFFFFFF0;
    // rom_array[40090] = 32'hFFFFFFF0;
    // rom_array[40091] = 32'hFFFFFFF1;
    // rom_array[40092] = 32'hFFFFFFF1;
    // rom_array[40093] = 32'hFFFFFFF0;
    // rom_array[40094] = 32'hFFFFFFF0;
    // rom_array[40095] = 32'hFFFFFFF0;
    // rom_array[40096] = 32'hFFFFFFF0;
    // rom_array[40097] = 32'hFFFFFFF0;
    // rom_array[40098] = 32'hFFFFFFF0;
    // rom_array[40099] = 32'hFFFFFFF1;
    // rom_array[40100] = 32'hFFFFFFF1;
    // rom_array[40101] = 32'hFFFFFFF0;
    // rom_array[40102] = 32'hFFFFFFF0;
    // rom_array[40103] = 32'hFFFFFFF0;
    // rom_array[40104] = 32'hFFFFFFF0;
    // rom_array[40105] = 32'hFFFFFFF1;
    // rom_array[40106] = 32'hFFFFFFF1;
    // rom_array[40107] = 32'hFFFFFFF1;
    // rom_array[40108] = 32'hFFFFFFF1;
    // rom_array[40109] = 32'hFFFFFFF1;
    // rom_array[40110] = 32'hFFFFFFF1;
    // rom_array[40111] = 32'hFFFFFFF1;
    // rom_array[40112] = 32'hFFFFFFF1;
    // rom_array[40113] = 32'hFFFFFFF1;
    // rom_array[40114] = 32'hFFFFFFF1;
    // rom_array[40115] = 32'hFFFFFFF1;
    // rom_array[40116] = 32'hFFFFFFF1;
    // rom_array[40117] = 32'hFFFFFFF1;
    // rom_array[40118] = 32'hFFFFFFF1;
    // rom_array[40119] = 32'hFFFFFFF1;
    // rom_array[40120] = 32'hFFFFFFF1;
    // rom_array[40121] = 32'hFFFFFFF1;
    // rom_array[40122] = 32'hFFFFFFF1;
    // rom_array[40123] = 32'hFFFFFFF1;
    // rom_array[40124] = 32'hFFFFFFF1;
    // rom_array[40125] = 32'hFFFFFFF1;
    // rom_array[40126] = 32'hFFFFFFF1;
    // rom_array[40127] = 32'hFFFFFFF1;
    // rom_array[40128] = 32'hFFFFFFF1;
    // rom_array[40129] = 32'hFFFFFFF1;
    // rom_array[40130] = 32'hFFFFFFF1;
    // rom_array[40131] = 32'hFFFFFFF1;
    // rom_array[40132] = 32'hFFFFFFF1;
    // rom_array[40133] = 32'hFFFFFFF1;
    // rom_array[40134] = 32'hFFFFFFF1;
    // rom_array[40135] = 32'hFFFFFFF1;
    // rom_array[40136] = 32'hFFFFFFF1;
    // rom_array[40137] = 32'hFFFFFFF1;
    // rom_array[40138] = 32'hFFFFFFF1;
    // rom_array[40139] = 32'hFFFFFFF1;
    // rom_array[40140] = 32'hFFFFFFF1;
    // rom_array[40141] = 32'hFFFFFFF1;
    // rom_array[40142] = 32'hFFFFFFF1;
    // rom_array[40143] = 32'hFFFFFFF1;
    // rom_array[40144] = 32'hFFFFFFF1;
    // rom_array[40145] = 32'hFFFFFFF1;
    // rom_array[40146] = 32'hFFFFFFF1;
    // rom_array[40147] = 32'hFFFFFFF1;
    // rom_array[40148] = 32'hFFFFFFF1;
    // rom_array[40149] = 32'hFFFFFFF1;
    // rom_array[40150] = 32'hFFFFFFF1;
    // rom_array[40151] = 32'hFFFFFFF1;
    // rom_array[40152] = 32'hFFFFFFF1;
    // rom_array[40153] = 32'hFFFFFFF1;
    // rom_array[40154] = 32'hFFFFFFF1;
    // rom_array[40155] = 32'hFFFFFFF1;
    // rom_array[40156] = 32'hFFFFFFF1;
    // rom_array[40157] = 32'hFFFFFFF1;
    // rom_array[40158] = 32'hFFFFFFF1;
    // rom_array[40159] = 32'hFFFFFFF1;
    // rom_array[40160] = 32'hFFFFFFF1;
    // rom_array[40161] = 32'hFFFFFFF1;
    // rom_array[40162] = 32'hFFFFFFF1;
    // rom_array[40163] = 32'hFFFFFFF1;
    // rom_array[40164] = 32'hFFFFFFF1;
    // rom_array[40165] = 32'hFFFFFFF1;
    // rom_array[40166] = 32'hFFFFFFF1;
    // rom_array[40167] = 32'hFFFFFFF1;
    // rom_array[40168] = 32'hFFFFFFF1;
    // rom_array[40169] = 32'hFFFFFFF1;
    // rom_array[40170] = 32'hFFFFFFF1;
    // rom_array[40171] = 32'hFFFFFFF1;
    // rom_array[40172] = 32'hFFFFFFF1;
    // rom_array[40173] = 32'hFFFFFFF1;
    // rom_array[40174] = 32'hFFFFFFF1;
    // rom_array[40175] = 32'hFFFFFFF1;
    // rom_array[40176] = 32'hFFFFFFF1;
    // rom_array[40177] = 32'hFFFFFFF1;
    // rom_array[40178] = 32'hFFFFFFF1;
    // rom_array[40179] = 32'hFFFFFFF1;
    // rom_array[40180] = 32'hFFFFFFF1;
    // rom_array[40181] = 32'hFFFFFFF1;
    // rom_array[40182] = 32'hFFFFFFF1;
    // rom_array[40183] = 32'hFFFFFFF1;
    // rom_array[40184] = 32'hFFFFFFF1;
    // rom_array[40185] = 32'hFFFFFFF1;
    // rom_array[40186] = 32'hFFFFFFF1;
    // rom_array[40187] = 32'hFFFFFFF1;
    // rom_array[40188] = 32'hFFFFFFF1;
    // rom_array[40189] = 32'hFFFFFFF1;
    // rom_array[40190] = 32'hFFFFFFF1;
    // rom_array[40191] = 32'hFFFFFFF1;
    // rom_array[40192] = 32'hFFFFFFF1;
    // rom_array[40193] = 32'hFFFFFFF1;
    // rom_array[40194] = 32'hFFFFFFF1;
    // rom_array[40195] = 32'hFFFFFFF1;
    // rom_array[40196] = 32'hFFFFFFF1;
    // rom_array[40197] = 32'hFFFFFFF1;
    // rom_array[40198] = 32'hFFFFFFF1;
    // rom_array[40199] = 32'hFFFFFFF1;
    // rom_array[40200] = 32'hFFFFFFF1;
    // rom_array[40201] = 32'hFFFFFFF1;
    // rom_array[40202] = 32'hFFFFFFF1;
    // rom_array[40203] = 32'hFFFFFFF1;
    // rom_array[40204] = 32'hFFFFFFF1;
    // rom_array[40205] = 32'hFFFFFFF1;
    // rom_array[40206] = 32'hFFFFFFF1;
    // rom_array[40207] = 32'hFFFFFFF1;
    // rom_array[40208] = 32'hFFFFFFF1;
    // rom_array[40209] = 32'hFFFFFFF1;
    // rom_array[40210] = 32'hFFFFFFF1;
    // rom_array[40211] = 32'hFFFFFFF1;
    // rom_array[40212] = 32'hFFFFFFF1;
    // rom_array[40213] = 32'hFFFFFFF1;
    // rom_array[40214] = 32'hFFFFFFF1;
    // rom_array[40215] = 32'hFFFFFFF1;
    // rom_array[40216] = 32'hFFFFFFF1;
    // rom_array[40217] = 32'hFFFFFFF1;
    // rom_array[40218] = 32'hFFFFFFF1;
    // rom_array[40219] = 32'hFFFFFFF1;
    // rom_array[40220] = 32'hFFFFFFF1;
    // rom_array[40221] = 32'hFFFFFFF1;
    // rom_array[40222] = 32'hFFFFFFF1;
    // rom_array[40223] = 32'hFFFFFFF1;
    // rom_array[40224] = 32'hFFFFFFF1;
    // rom_array[40225] = 32'hFFFFFFF1;
    // rom_array[40226] = 32'hFFFFFFF1;
    // rom_array[40227] = 32'hFFFFFFF1;
    // rom_array[40228] = 32'hFFFFFFF1;
    // rom_array[40229] = 32'hFFFFFFF1;
    // rom_array[40230] = 32'hFFFFFFF1;
    // rom_array[40231] = 32'hFFFFFFF1;
    // rom_array[40232] = 32'hFFFFFFF1;
    // rom_array[40233] = 32'hFFFFFFF1;
    // rom_array[40234] = 32'hFFFFFFF1;
    // rom_array[40235] = 32'hFFFFFFF1;
    // rom_array[40236] = 32'hFFFFFFF1;
    // rom_array[40237] = 32'hFFFFFFF0;
    // rom_array[40238] = 32'hFFFFFFF0;
    // rom_array[40239] = 32'hFFFFFFF0;
    // rom_array[40240] = 32'hFFFFFFF0;
    // rom_array[40241] = 32'hFFFFFFF1;
    // rom_array[40242] = 32'hFFFFFFF1;
    // rom_array[40243] = 32'hFFFFFFF1;
    // rom_array[40244] = 32'hFFFFFFF1;
    // rom_array[40245] = 32'hFFFFFFF0;
    // rom_array[40246] = 32'hFFFFFFF0;
    // rom_array[40247] = 32'hFFFFFFF0;
    // rom_array[40248] = 32'hFFFFFFF0;
    // rom_array[40249] = 32'hFFFFFFF1;
    // rom_array[40250] = 32'hFFFFFFF1;
    // rom_array[40251] = 32'hFFFFFFF1;
    // rom_array[40252] = 32'hFFFFFFF1;
    // rom_array[40253] = 32'hFFFFFFF0;
    // rom_array[40254] = 32'hFFFFFFF0;
    // rom_array[40255] = 32'hFFFFFFF0;
    // rom_array[40256] = 32'hFFFFFFF0;
    // rom_array[40257] = 32'hFFFFFFF1;
    // rom_array[40258] = 32'hFFFFFFF1;
    // rom_array[40259] = 32'hFFFFFFF1;
    // rom_array[40260] = 32'hFFFFFFF1;
    // rom_array[40261] = 32'hFFFFFFF0;
    // rom_array[40262] = 32'hFFFFFFF0;
    // rom_array[40263] = 32'hFFFFFFF0;
    // rom_array[40264] = 32'hFFFFFFF0;
    // rom_array[40265] = 32'hFFFFFFF1;
    // rom_array[40266] = 32'hFFFFFFF1;
    // rom_array[40267] = 32'hFFFFFFF1;
    // rom_array[40268] = 32'hFFFFFFF1;
    // rom_array[40269] = 32'hFFFFFFF0;
    // rom_array[40270] = 32'hFFFFFFF0;
    // rom_array[40271] = 32'hFFFFFFF0;
    // rom_array[40272] = 32'hFFFFFFF0;
    // rom_array[40273] = 32'hFFFFFFF1;
    // rom_array[40274] = 32'hFFFFFFF1;
    // rom_array[40275] = 32'hFFFFFFF1;
    // rom_array[40276] = 32'hFFFFFFF1;
    // rom_array[40277] = 32'hFFFFFFF0;
    // rom_array[40278] = 32'hFFFFFFF0;
    // rom_array[40279] = 32'hFFFFFFF0;
    // rom_array[40280] = 32'hFFFFFFF0;
    // rom_array[40281] = 32'hFFFFFFF1;
    // rom_array[40282] = 32'hFFFFFFF1;
    // rom_array[40283] = 32'hFFFFFFF1;
    // rom_array[40284] = 32'hFFFFFFF1;
    // rom_array[40285] = 32'hFFFFFFF0;
    // rom_array[40286] = 32'hFFFFFFF0;
    // rom_array[40287] = 32'hFFFFFFF0;
    // rom_array[40288] = 32'hFFFFFFF0;
    // rom_array[40289] = 32'hFFFFFFF1;
    // rom_array[40290] = 32'hFFFFFFF1;
    // rom_array[40291] = 32'hFFFFFFF1;
    // rom_array[40292] = 32'hFFFFFFF1;
    // rom_array[40293] = 32'hFFFFFFF0;
    // rom_array[40294] = 32'hFFFFFFF0;
    // rom_array[40295] = 32'hFFFFFFF0;
    // rom_array[40296] = 32'hFFFFFFF0;
    // rom_array[40297] = 32'hFFFFFFF1;
    // rom_array[40298] = 32'hFFFFFFF1;
    // rom_array[40299] = 32'hFFFFFFF1;
    // rom_array[40300] = 32'hFFFFFFF1;
    // rom_array[40301] = 32'hFFFFFFF0;
    // rom_array[40302] = 32'hFFFFFFF0;
    // rom_array[40303] = 32'hFFFFFFF0;
    // rom_array[40304] = 32'hFFFFFFF0;
    // rom_array[40305] = 32'hFFFFFFF1;
    // rom_array[40306] = 32'hFFFFFFF1;
    // rom_array[40307] = 32'hFFFFFFF1;
    // rom_array[40308] = 32'hFFFFFFF1;
    // rom_array[40309] = 32'hFFFFFFF0;
    // rom_array[40310] = 32'hFFFFFFF0;
    // rom_array[40311] = 32'hFFFFFFF0;
    // rom_array[40312] = 32'hFFFFFFF0;
    // rom_array[40313] = 32'hFFFFFFF1;
    // rom_array[40314] = 32'hFFFFFFF1;
    // rom_array[40315] = 32'hFFFFFFF1;
    // rom_array[40316] = 32'hFFFFFFF1;
    // rom_array[40317] = 32'hFFFFFFF0;
    // rom_array[40318] = 32'hFFFFFFF0;
    // rom_array[40319] = 32'hFFFFFFF0;
    // rom_array[40320] = 32'hFFFFFFF0;
    // rom_array[40321] = 32'hFFFFFFF1;
    // rom_array[40322] = 32'hFFFFFFF1;
    // rom_array[40323] = 32'hFFFFFFF1;
    // rom_array[40324] = 32'hFFFFFFF1;
    // rom_array[40325] = 32'hFFFFFFF0;
    // rom_array[40326] = 32'hFFFFFFF0;
    // rom_array[40327] = 32'hFFFFFFF0;
    // rom_array[40328] = 32'hFFFFFFF0;
    // rom_array[40329] = 32'hFFFFFFF1;
    // rom_array[40330] = 32'hFFFFFFF1;
    // rom_array[40331] = 32'hFFFFFFF1;
    // rom_array[40332] = 32'hFFFFFFF1;
    // rom_array[40333] = 32'hFFFFFFF0;
    // rom_array[40334] = 32'hFFFFFFF0;
    // rom_array[40335] = 32'hFFFFFFF0;
    // rom_array[40336] = 32'hFFFFFFF0;
    // rom_array[40337] = 32'hFFFFFFF1;
    // rom_array[40338] = 32'hFFFFFFF1;
    // rom_array[40339] = 32'hFFFFFFF1;
    // rom_array[40340] = 32'hFFFFFFF1;
    // rom_array[40341] = 32'hFFFFFFF0;
    // rom_array[40342] = 32'hFFFFFFF0;
    // rom_array[40343] = 32'hFFFFFFF0;
    // rom_array[40344] = 32'hFFFFFFF0;
    // rom_array[40345] = 32'hFFFFFFF1;
    // rom_array[40346] = 32'hFFFFFFF1;
    // rom_array[40347] = 32'hFFFFFFF1;
    // rom_array[40348] = 32'hFFFFFFF1;
    // rom_array[40349] = 32'hFFFFFFF0;
    // rom_array[40350] = 32'hFFFFFFF0;
    // rom_array[40351] = 32'hFFFFFFF0;
    // rom_array[40352] = 32'hFFFFFFF0;
    // rom_array[40353] = 32'hFFFFFFF1;
    // rom_array[40354] = 32'hFFFFFFF1;
    // rom_array[40355] = 32'hFFFFFFF1;
    // rom_array[40356] = 32'hFFFFFFF1;
    // rom_array[40357] = 32'hFFFFFFF0;
    // rom_array[40358] = 32'hFFFFFFF0;
    // rom_array[40359] = 32'hFFFFFFF0;
    // rom_array[40360] = 32'hFFFFFFF0;
    // rom_array[40361] = 32'hFFFFFFF1;
    // rom_array[40362] = 32'hFFFFFFF1;
    // rom_array[40363] = 32'hFFFFFFF1;
    // rom_array[40364] = 32'hFFFFFFF1;
    // rom_array[40365] = 32'hFFFFFFF0;
    // rom_array[40366] = 32'hFFFFFFF0;
    // rom_array[40367] = 32'hFFFFFFF0;
    // rom_array[40368] = 32'hFFFFFFF0;
    // rom_array[40369] = 32'hFFFFFFF1;
    // rom_array[40370] = 32'hFFFFFFF1;
    // rom_array[40371] = 32'hFFFFFFF1;
    // rom_array[40372] = 32'hFFFFFFF1;
    // rom_array[40373] = 32'hFFFFFFF0;
    // rom_array[40374] = 32'hFFFFFFF0;
    // rom_array[40375] = 32'hFFFFFFF0;
    // rom_array[40376] = 32'hFFFFFFF0;
    // rom_array[40377] = 32'hFFFFFFF1;
    // rom_array[40378] = 32'hFFFFFFF1;
    // rom_array[40379] = 32'hFFFFFFF1;
    // rom_array[40380] = 32'hFFFFFFF1;
    // rom_array[40381] = 32'hFFFFFFF1;
    // rom_array[40382] = 32'hFFFFFFF1;
    // rom_array[40383] = 32'hFFFFFFF1;
    // rom_array[40384] = 32'hFFFFFFF1;
    // rom_array[40385] = 32'hFFFFFFF1;
    // rom_array[40386] = 32'hFFFFFFF1;
    // rom_array[40387] = 32'hFFFFFFF1;
    // rom_array[40388] = 32'hFFFFFFF1;
    // rom_array[40389] = 32'hFFFFFFF1;
    // rom_array[40390] = 32'hFFFFFFF1;
    // rom_array[40391] = 32'hFFFFFFF1;
    // rom_array[40392] = 32'hFFFFFFF1;
    // rom_array[40393] = 32'hFFFFFFF1;
    // rom_array[40394] = 32'hFFFFFFF1;
    // rom_array[40395] = 32'hFFFFFFF1;
    // rom_array[40396] = 32'hFFFFFFF1;
    // rom_array[40397] = 32'hFFFFFFF0;
    // rom_array[40398] = 32'hFFFFFFF0;
    // rom_array[40399] = 32'hFFFFFFF0;
    // rom_array[40400] = 32'hFFFFFFF0;
    // rom_array[40401] = 32'hFFFFFFF1;
    // rom_array[40402] = 32'hFFFFFFF1;
    // rom_array[40403] = 32'hFFFFFFF1;
    // rom_array[40404] = 32'hFFFFFFF1;
    // rom_array[40405] = 32'hFFFFFFF0;
    // rom_array[40406] = 32'hFFFFFFF0;
    // rom_array[40407] = 32'hFFFFFFF0;
    // rom_array[40408] = 32'hFFFFFFF0;
    // rom_array[40409] = 32'hFFFFFFF1;
    // rom_array[40410] = 32'hFFFFFFF1;
    // rom_array[40411] = 32'hFFFFFFF1;
    // rom_array[40412] = 32'hFFFFFFF1;
    // rom_array[40413] = 32'hFFFFFFF0;
    // rom_array[40414] = 32'hFFFFFFF0;
    // rom_array[40415] = 32'hFFFFFFF0;
    // rom_array[40416] = 32'hFFFFFFF0;
    // rom_array[40417] = 32'hFFFFFFF1;
    // rom_array[40418] = 32'hFFFFFFF1;
    // rom_array[40419] = 32'hFFFFFFF1;
    // rom_array[40420] = 32'hFFFFFFF1;
    // rom_array[40421] = 32'hFFFFFFF0;
    // rom_array[40422] = 32'hFFFFFFF0;
    // rom_array[40423] = 32'hFFFFFFF0;
    // rom_array[40424] = 32'hFFFFFFF0;
    // rom_array[40425] = 32'hFFFFFFF0;
    // rom_array[40426] = 32'hFFFFFFF0;
    // rom_array[40427] = 32'hFFFFFFF0;
    // rom_array[40428] = 32'hFFFFFFF0;
    // rom_array[40429] = 32'hFFFFFFF0;
    // rom_array[40430] = 32'hFFFFFFF0;
    // rom_array[40431] = 32'hFFFFFFF1;
    // rom_array[40432] = 32'hFFFFFFF1;
    // rom_array[40433] = 32'hFFFFFFF0;
    // rom_array[40434] = 32'hFFFFFFF0;
    // rom_array[40435] = 32'hFFFFFFF0;
    // rom_array[40436] = 32'hFFFFFFF0;
    // rom_array[40437] = 32'hFFFFFFF0;
    // rom_array[40438] = 32'hFFFFFFF0;
    // rom_array[40439] = 32'hFFFFFFF1;
    // rom_array[40440] = 32'hFFFFFFF1;
    // rom_array[40441] = 32'hFFFFFFF0;
    // rom_array[40442] = 32'hFFFFFFF0;
    // rom_array[40443] = 32'hFFFFFFF0;
    // rom_array[40444] = 32'hFFFFFFF0;
    // rom_array[40445] = 32'hFFFFFFF1;
    // rom_array[40446] = 32'hFFFFFFF1;
    // rom_array[40447] = 32'hFFFFFFF1;
    // rom_array[40448] = 32'hFFFFFFF1;
    // rom_array[40449] = 32'hFFFFFFF0;
    // rom_array[40450] = 32'hFFFFFFF0;
    // rom_array[40451] = 32'hFFFFFFF0;
    // rom_array[40452] = 32'hFFFFFFF0;
    // rom_array[40453] = 32'hFFFFFFF1;
    // rom_array[40454] = 32'hFFFFFFF1;
    // rom_array[40455] = 32'hFFFFFFF1;
    // rom_array[40456] = 32'hFFFFFFF1;
    // rom_array[40457] = 32'hFFFFFFF0;
    // rom_array[40458] = 32'hFFFFFFF0;
    // rom_array[40459] = 32'hFFFFFFF1;
    // rom_array[40460] = 32'hFFFFFFF1;
    // rom_array[40461] = 32'hFFFFFFF0;
    // rom_array[40462] = 32'hFFFFFFF0;
    // rom_array[40463] = 32'hFFFFFFF1;
    // rom_array[40464] = 32'hFFFFFFF1;
    // rom_array[40465] = 32'hFFFFFFF0;
    // rom_array[40466] = 32'hFFFFFFF0;
    // rom_array[40467] = 32'hFFFFFFF1;
    // rom_array[40468] = 32'hFFFFFFF1;
    // rom_array[40469] = 32'hFFFFFFF0;
    // rom_array[40470] = 32'hFFFFFFF0;
    // rom_array[40471] = 32'hFFFFFFF1;
    // rom_array[40472] = 32'hFFFFFFF1;
    // rom_array[40473] = 32'hFFFFFFF0;
    // rom_array[40474] = 32'hFFFFFFF0;
    // rom_array[40475] = 32'hFFFFFFF1;
    // rom_array[40476] = 32'hFFFFFFF1;
    // rom_array[40477] = 32'hFFFFFFF0;
    // rom_array[40478] = 32'hFFFFFFF0;
    // rom_array[40479] = 32'hFFFFFFF1;
    // rom_array[40480] = 32'hFFFFFFF1;
    // rom_array[40481] = 32'hFFFFFFF0;
    // rom_array[40482] = 32'hFFFFFFF0;
    // rom_array[40483] = 32'hFFFFFFF1;
    // rom_array[40484] = 32'hFFFFFFF1;
    // rom_array[40485] = 32'hFFFFFFF0;
    // rom_array[40486] = 32'hFFFFFFF0;
    // rom_array[40487] = 32'hFFFFFFF1;
    // rom_array[40488] = 32'hFFFFFFF1;
    // rom_array[40489] = 32'hFFFFFFF0;
    // rom_array[40490] = 32'hFFFFFFF0;
    // rom_array[40491] = 32'hFFFFFFF0;
    // rom_array[40492] = 32'hFFFFFFF0;
    // rom_array[40493] = 32'hFFFFFFF1;
    // rom_array[40494] = 32'hFFFFFFF1;
    // rom_array[40495] = 32'hFFFFFFF1;
    // rom_array[40496] = 32'hFFFFFFF1;
    // rom_array[40497] = 32'hFFFFFFF0;
    // rom_array[40498] = 32'hFFFFFFF0;
    // rom_array[40499] = 32'hFFFFFFF0;
    // rom_array[40500] = 32'hFFFFFFF0;
    // rom_array[40501] = 32'hFFFFFFF1;
    // rom_array[40502] = 32'hFFFFFFF1;
    // rom_array[40503] = 32'hFFFFFFF1;
    // rom_array[40504] = 32'hFFFFFFF1;
    // rom_array[40505] = 32'hFFFFFFF0;
    // rom_array[40506] = 32'hFFFFFFF0;
    // rom_array[40507] = 32'hFFFFFFF0;
    // rom_array[40508] = 32'hFFFFFFF0;
    // rom_array[40509] = 32'hFFFFFFF1;
    // rom_array[40510] = 32'hFFFFFFF1;
    // rom_array[40511] = 32'hFFFFFFF1;
    // rom_array[40512] = 32'hFFFFFFF1;
    // rom_array[40513] = 32'hFFFFFFF0;
    // rom_array[40514] = 32'hFFFFFFF0;
    // rom_array[40515] = 32'hFFFFFFF0;
    // rom_array[40516] = 32'hFFFFFFF0;
    // rom_array[40517] = 32'hFFFFFFF1;
    // rom_array[40518] = 32'hFFFFFFF1;
    // rom_array[40519] = 32'hFFFFFFF1;
    // rom_array[40520] = 32'hFFFFFFF1;
    // rom_array[40521] = 32'hFFFFFFF0;
    // rom_array[40522] = 32'hFFFFFFF0;
    // rom_array[40523] = 32'hFFFFFFF0;
    // rom_array[40524] = 32'hFFFFFFF0;
    // rom_array[40525] = 32'hFFFFFFF1;
    // rom_array[40526] = 32'hFFFFFFF1;
    // rom_array[40527] = 32'hFFFFFFF1;
    // rom_array[40528] = 32'hFFFFFFF1;
    // rom_array[40529] = 32'hFFFFFFF0;
    // rom_array[40530] = 32'hFFFFFFF0;
    // rom_array[40531] = 32'hFFFFFFF0;
    // rom_array[40532] = 32'hFFFFFFF0;
    // rom_array[40533] = 32'hFFFFFFF1;
    // rom_array[40534] = 32'hFFFFFFF1;
    // rom_array[40535] = 32'hFFFFFFF1;
    // rom_array[40536] = 32'hFFFFFFF1;
    // rom_array[40537] = 32'hFFFFFFF0;
    // rom_array[40538] = 32'hFFFFFFF0;
    // rom_array[40539] = 32'hFFFFFFF0;
    // rom_array[40540] = 32'hFFFFFFF0;
    // rom_array[40541] = 32'hFFFFFFF1;
    // rom_array[40542] = 32'hFFFFFFF1;
    // rom_array[40543] = 32'hFFFFFFF1;
    // rom_array[40544] = 32'hFFFFFFF1;
    // rom_array[40545] = 32'hFFFFFFF0;
    // rom_array[40546] = 32'hFFFFFFF0;
    // rom_array[40547] = 32'hFFFFFFF0;
    // rom_array[40548] = 32'hFFFFFFF0;
    // rom_array[40549] = 32'hFFFFFFF1;
    // rom_array[40550] = 32'hFFFFFFF1;
    // rom_array[40551] = 32'hFFFFFFF1;
    // rom_array[40552] = 32'hFFFFFFF1;
    // rom_array[40553] = 32'hFFFFFFF0;
    // rom_array[40554] = 32'hFFFFFFF0;
    // rom_array[40555] = 32'hFFFFFFF1;
    // rom_array[40556] = 32'hFFFFFFF1;
    // rom_array[40557] = 32'hFFFFFFF0;
    // rom_array[40558] = 32'hFFFFFFF0;
    // rom_array[40559] = 32'hFFFFFFF1;
    // rom_array[40560] = 32'hFFFFFFF1;
    // rom_array[40561] = 32'hFFFFFFF0;
    // rom_array[40562] = 32'hFFFFFFF0;
    // rom_array[40563] = 32'hFFFFFFF1;
    // rom_array[40564] = 32'hFFFFFFF1;
    // rom_array[40565] = 32'hFFFFFFF0;
    // rom_array[40566] = 32'hFFFFFFF0;
    // rom_array[40567] = 32'hFFFFFFF1;
    // rom_array[40568] = 32'hFFFFFFF1;
    // rom_array[40569] = 32'hFFFFFFF0;
    // rom_array[40570] = 32'hFFFFFFF0;
    // rom_array[40571] = 32'hFFFFFFF1;
    // rom_array[40572] = 32'hFFFFFFF1;
    // rom_array[40573] = 32'hFFFFFFF0;
    // rom_array[40574] = 32'hFFFFFFF0;
    // rom_array[40575] = 32'hFFFFFFF1;
    // rom_array[40576] = 32'hFFFFFFF1;
    // rom_array[40577] = 32'hFFFFFFF0;
    // rom_array[40578] = 32'hFFFFFFF0;
    // rom_array[40579] = 32'hFFFFFFF1;
    // rom_array[40580] = 32'hFFFFFFF1;
    // rom_array[40581] = 32'hFFFFFFF0;
    // rom_array[40582] = 32'hFFFFFFF0;
    // rom_array[40583] = 32'hFFFFFFF1;
    // rom_array[40584] = 32'hFFFFFFF1;
    // rom_array[40585] = 32'hFFFFFFF0;
    // rom_array[40586] = 32'hFFFFFFF0;
    // rom_array[40587] = 32'hFFFFFFF0;
    // rom_array[40588] = 32'hFFFFFFF0;
    // rom_array[40589] = 32'hFFFFFFF1;
    // rom_array[40590] = 32'hFFFFFFF1;
    // rom_array[40591] = 32'hFFFFFFF1;
    // rom_array[40592] = 32'hFFFFFFF1;
    // rom_array[40593] = 32'hFFFFFFF0;
    // rom_array[40594] = 32'hFFFFFFF0;
    // rom_array[40595] = 32'hFFFFFFF0;
    // rom_array[40596] = 32'hFFFFFFF0;
    // rom_array[40597] = 32'hFFFFFFF1;
    // rom_array[40598] = 32'hFFFFFFF1;
    // rom_array[40599] = 32'hFFFFFFF1;
    // rom_array[40600] = 32'hFFFFFFF1;
    // rom_array[40601] = 32'hFFFFFFF0;
    // rom_array[40602] = 32'hFFFFFFF0;
    // rom_array[40603] = 32'hFFFFFFF0;
    // rom_array[40604] = 32'hFFFFFFF0;
    // rom_array[40605] = 32'hFFFFFFF1;
    // rom_array[40606] = 32'hFFFFFFF1;
    // rom_array[40607] = 32'hFFFFFFF1;
    // rom_array[40608] = 32'hFFFFFFF1;
    // rom_array[40609] = 32'hFFFFFFF0;
    // rom_array[40610] = 32'hFFFFFFF0;
    // rom_array[40611] = 32'hFFFFFFF0;
    // rom_array[40612] = 32'hFFFFFFF0;
    // rom_array[40613] = 32'hFFFFFFF1;
    // rom_array[40614] = 32'hFFFFFFF1;
    // rom_array[40615] = 32'hFFFFFFF1;
    // rom_array[40616] = 32'hFFFFFFF1;
    // rom_array[40617] = 32'hFFFFFFF0;
    // rom_array[40618] = 32'hFFFFFFF0;
    // rom_array[40619] = 32'hFFFFFFF1;
    // rom_array[40620] = 32'hFFFFFFF1;
    // rom_array[40621] = 32'hFFFFFFF1;
    // rom_array[40622] = 32'hFFFFFFF1;
    // rom_array[40623] = 32'hFFFFFFF1;
    // rom_array[40624] = 32'hFFFFFFF1;
    // rom_array[40625] = 32'hFFFFFFF0;
    // rom_array[40626] = 32'hFFFFFFF0;
    // rom_array[40627] = 32'hFFFFFFF1;
    // rom_array[40628] = 32'hFFFFFFF1;
    // rom_array[40629] = 32'hFFFFFFF1;
    // rom_array[40630] = 32'hFFFFFFF1;
    // rom_array[40631] = 32'hFFFFFFF1;
    // rom_array[40632] = 32'hFFFFFFF1;
    // rom_array[40633] = 32'hFFFFFFF1;
    // rom_array[40634] = 32'hFFFFFFF1;
    // rom_array[40635] = 32'hFFFFFFF1;
    // rom_array[40636] = 32'hFFFFFFF1;
    // rom_array[40637] = 32'hFFFFFFF1;
    // rom_array[40638] = 32'hFFFFFFF1;
    // rom_array[40639] = 32'hFFFFFFF1;
    // rom_array[40640] = 32'hFFFFFFF1;
    // rom_array[40641] = 32'hFFFFFFF1;
    // rom_array[40642] = 32'hFFFFFFF1;
    // rom_array[40643] = 32'hFFFFFFF1;
    // rom_array[40644] = 32'hFFFFFFF1;
    // rom_array[40645] = 32'hFFFFFFF1;
    // rom_array[40646] = 32'hFFFFFFF1;
    // rom_array[40647] = 32'hFFFFFFF1;
    // rom_array[40648] = 32'hFFFFFFF1;
    // rom_array[40649] = 32'hFFFFFFF0;
    // rom_array[40650] = 32'hFFFFFFF0;
    // rom_array[40651] = 32'hFFFFFFF0;
    // rom_array[40652] = 32'hFFFFFFF0;
    // rom_array[40653] = 32'hFFFFFFF1;
    // rom_array[40654] = 32'hFFFFFFF1;
    // rom_array[40655] = 32'hFFFFFFF1;
    // rom_array[40656] = 32'hFFFFFFF1;
    // rom_array[40657] = 32'hFFFFFFF0;
    // rom_array[40658] = 32'hFFFFFFF0;
    // rom_array[40659] = 32'hFFFFFFF0;
    // rom_array[40660] = 32'hFFFFFFF0;
    // rom_array[40661] = 32'hFFFFFFF1;
    // rom_array[40662] = 32'hFFFFFFF1;
    // rom_array[40663] = 32'hFFFFFFF1;
    // rom_array[40664] = 32'hFFFFFFF1;
    // rom_array[40665] = 32'hFFFFFFF0;
    // rom_array[40666] = 32'hFFFFFFF0;
    // rom_array[40667] = 32'hFFFFFFF0;
    // rom_array[40668] = 32'hFFFFFFF0;
    // rom_array[40669] = 32'hFFFFFFF1;
    // rom_array[40670] = 32'hFFFFFFF1;
    // rom_array[40671] = 32'hFFFFFFF1;
    // rom_array[40672] = 32'hFFFFFFF1;
    // rom_array[40673] = 32'hFFFFFFF0;
    // rom_array[40674] = 32'hFFFFFFF0;
    // rom_array[40675] = 32'hFFFFFFF0;
    // rom_array[40676] = 32'hFFFFFFF0;
    // rom_array[40677] = 32'hFFFFFFF1;
    // rom_array[40678] = 32'hFFFFFFF1;
    // rom_array[40679] = 32'hFFFFFFF1;
    // rom_array[40680] = 32'hFFFFFFF1;
    // rom_array[40681] = 32'hFFFFFFF0;
    // rom_array[40682] = 32'hFFFFFFF0;
    // rom_array[40683] = 32'hFFFFFFF0;
    // rom_array[40684] = 32'hFFFFFFF0;
    // rom_array[40685] = 32'hFFFFFFF1;
    // rom_array[40686] = 32'hFFFFFFF1;
    // rom_array[40687] = 32'hFFFFFFF1;
    // rom_array[40688] = 32'hFFFFFFF1;
    // rom_array[40689] = 32'hFFFFFFF0;
    // rom_array[40690] = 32'hFFFFFFF0;
    // rom_array[40691] = 32'hFFFFFFF0;
    // rom_array[40692] = 32'hFFFFFFF0;
    // rom_array[40693] = 32'hFFFFFFF1;
    // rom_array[40694] = 32'hFFFFFFF1;
    // rom_array[40695] = 32'hFFFFFFF1;
    // rom_array[40696] = 32'hFFFFFFF1;
    // rom_array[40697] = 32'hFFFFFFF1;
    // rom_array[40698] = 32'hFFFFFFF1;
    // rom_array[40699] = 32'hFFFFFFF1;
    // rom_array[40700] = 32'hFFFFFFF1;
    // rom_array[40701] = 32'hFFFFFFF1;
    // rom_array[40702] = 32'hFFFFFFF1;
    // rom_array[40703] = 32'hFFFFFFF1;
    // rom_array[40704] = 32'hFFFFFFF1;
    // rom_array[40705] = 32'hFFFFFFF1;
    // rom_array[40706] = 32'hFFFFFFF1;
    // rom_array[40707] = 32'hFFFFFFF1;
    // rom_array[40708] = 32'hFFFFFFF1;
    // rom_array[40709] = 32'hFFFFFFF1;
    // rom_array[40710] = 32'hFFFFFFF1;
    // rom_array[40711] = 32'hFFFFFFF1;
    // rom_array[40712] = 32'hFFFFFFF1;
    // rom_array[40713] = 32'hFFFFFFF1;
    // rom_array[40714] = 32'hFFFFFFF1;
    // rom_array[40715] = 32'hFFFFFFF1;
    // rom_array[40716] = 32'hFFFFFFF1;
    // rom_array[40717] = 32'hFFFFFFF1;
    // rom_array[40718] = 32'hFFFFFFF1;
    // rom_array[40719] = 32'hFFFFFFF1;
    // rom_array[40720] = 32'hFFFFFFF1;
    // rom_array[40721] = 32'hFFFFFFF1;
    // rom_array[40722] = 32'hFFFFFFF1;
    // rom_array[40723] = 32'hFFFFFFF1;
    // rom_array[40724] = 32'hFFFFFFF1;
    // rom_array[40725] = 32'hFFFFFFF1;
    // rom_array[40726] = 32'hFFFFFFF1;
    // rom_array[40727] = 32'hFFFFFFF1;
    // rom_array[40728] = 32'hFFFFFFF1;
    // rom_array[40729] = 32'hFFFFFFF1;
    // rom_array[40730] = 32'hFFFFFFF1;
    // rom_array[40731] = 32'hFFFFFFF1;
    // rom_array[40732] = 32'hFFFFFFF1;
    // rom_array[40733] = 32'hFFFFFFF1;
    // rom_array[40734] = 32'hFFFFFFF1;
    // rom_array[40735] = 32'hFFFFFFF1;
    // rom_array[40736] = 32'hFFFFFFF1;
    // rom_array[40737] = 32'hFFFFFFF1;
    // rom_array[40738] = 32'hFFFFFFF1;
    // rom_array[40739] = 32'hFFFFFFF1;
    // rom_array[40740] = 32'hFFFFFFF1;
    // rom_array[40741] = 32'hFFFFFFF1;
    // rom_array[40742] = 32'hFFFFFFF1;
    // rom_array[40743] = 32'hFFFFFFF1;
    // rom_array[40744] = 32'hFFFFFFF1;
    // rom_array[40745] = 32'hFFFFFFF1;
    // rom_array[40746] = 32'hFFFFFFF1;
    // rom_array[40747] = 32'hFFFFFFF1;
    // rom_array[40748] = 32'hFFFFFFF1;
    // rom_array[40749] = 32'hFFFFFFF1;
    // rom_array[40750] = 32'hFFFFFFF1;
    // rom_array[40751] = 32'hFFFFFFF1;
    // rom_array[40752] = 32'hFFFFFFF1;
    // rom_array[40753] = 32'hFFFFFFF1;
    // rom_array[40754] = 32'hFFFFFFF1;
    // rom_array[40755] = 32'hFFFFFFF1;
    // rom_array[40756] = 32'hFFFFFFF1;
    // rom_array[40757] = 32'hFFFFFFF1;
    // rom_array[40758] = 32'hFFFFFFF1;
    // rom_array[40759] = 32'hFFFFFFF1;
    // rom_array[40760] = 32'hFFFFFFF1;
    // rom_array[40761] = 32'hFFFFFFF1;
    // rom_array[40762] = 32'hFFFFFFF1;
    // rom_array[40763] = 32'hFFFFFFF1;
    // rom_array[40764] = 32'hFFFFFFF1;
    // rom_array[40765] = 32'hFFFFFFF1;
    // rom_array[40766] = 32'hFFFFFFF1;
    // rom_array[40767] = 32'hFFFFFFF1;
    // rom_array[40768] = 32'hFFFFFFF1;
    // rom_array[40769] = 32'hFFFFFFF1;
    // rom_array[40770] = 32'hFFFFFFF1;
    // rom_array[40771] = 32'hFFFFFFF1;
    // rom_array[40772] = 32'hFFFFFFF1;
    // rom_array[40773] = 32'hFFFFFFF1;
    // rom_array[40774] = 32'hFFFFFFF1;
    // rom_array[40775] = 32'hFFFFFFF1;
    // rom_array[40776] = 32'hFFFFFFF1;
    // rom_array[40777] = 32'hFFFFFFF1;
    // rom_array[40778] = 32'hFFFFFFF1;
    // rom_array[40779] = 32'hFFFFFFF1;
    // rom_array[40780] = 32'hFFFFFFF1;
    // rom_array[40781] = 32'hFFFFFFF1;
    // rom_array[40782] = 32'hFFFFFFF1;
    // rom_array[40783] = 32'hFFFFFFF1;
    // rom_array[40784] = 32'hFFFFFFF1;
    // rom_array[40785] = 32'hFFFFFFF1;
    // rom_array[40786] = 32'hFFFFFFF1;
    // rom_array[40787] = 32'hFFFFFFF1;
    // rom_array[40788] = 32'hFFFFFFF1;
    // rom_array[40789] = 32'hFFFFFFF1;
    // rom_array[40790] = 32'hFFFFFFF1;
    // rom_array[40791] = 32'hFFFFFFF1;
    // rom_array[40792] = 32'hFFFFFFF1;
    // rom_array[40793] = 32'hFFFFFFF1;
    // rom_array[40794] = 32'hFFFFFFF1;
    // rom_array[40795] = 32'hFFFFFFF1;
    // rom_array[40796] = 32'hFFFFFFF1;
    // rom_array[40797] = 32'hFFFFFFF0;
    // rom_array[40798] = 32'hFFFFFFF0;
    // rom_array[40799] = 32'hFFFFFFF0;
    // rom_array[40800] = 32'hFFFFFFF0;
    // rom_array[40801] = 32'hFFFFFFF1;
    // rom_array[40802] = 32'hFFFFFFF1;
    // rom_array[40803] = 32'hFFFFFFF1;
    // rom_array[40804] = 32'hFFFFFFF1;
    // rom_array[40805] = 32'hFFFFFFF0;
    // rom_array[40806] = 32'hFFFFFFF0;
    // rom_array[40807] = 32'hFFFFFFF0;
    // rom_array[40808] = 32'hFFFFFFF0;
    // rom_array[40809] = 32'hFFFFFFF1;
    // rom_array[40810] = 32'hFFFFFFF1;
    // rom_array[40811] = 32'hFFFFFFF1;
    // rom_array[40812] = 32'hFFFFFFF1;
    // rom_array[40813] = 32'hFFFFFFF0;
    // rom_array[40814] = 32'hFFFFFFF0;
    // rom_array[40815] = 32'hFFFFFFF0;
    // rom_array[40816] = 32'hFFFFFFF0;
    // rom_array[40817] = 32'hFFFFFFF1;
    // rom_array[40818] = 32'hFFFFFFF1;
    // rom_array[40819] = 32'hFFFFFFF1;
    // rom_array[40820] = 32'hFFFFFFF1;
    // rom_array[40821] = 32'hFFFFFFF0;
    // rom_array[40822] = 32'hFFFFFFF0;
    // rom_array[40823] = 32'hFFFFFFF0;
    // rom_array[40824] = 32'hFFFFFFF0;
    // rom_array[40825] = 32'hFFFFFFF1;
    // rom_array[40826] = 32'hFFFFFFF1;
    // rom_array[40827] = 32'hFFFFFFF1;
    // rom_array[40828] = 32'hFFFFFFF1;
    // rom_array[40829] = 32'hFFFFFFF0;
    // rom_array[40830] = 32'hFFFFFFF0;
    // rom_array[40831] = 32'hFFFFFFF0;
    // rom_array[40832] = 32'hFFFFFFF0;
    // rom_array[40833] = 32'hFFFFFFF1;
    // rom_array[40834] = 32'hFFFFFFF1;
    // rom_array[40835] = 32'hFFFFFFF1;
    // rom_array[40836] = 32'hFFFFFFF1;
    // rom_array[40837] = 32'hFFFFFFF0;
    // rom_array[40838] = 32'hFFFFFFF0;
    // rom_array[40839] = 32'hFFFFFFF0;
    // rom_array[40840] = 32'hFFFFFFF0;
    // rom_array[40841] = 32'hFFFFFFF1;
    // rom_array[40842] = 32'hFFFFFFF1;
    // rom_array[40843] = 32'hFFFFFFF1;
    // rom_array[40844] = 32'hFFFFFFF1;
    // rom_array[40845] = 32'hFFFFFFF0;
    // rom_array[40846] = 32'hFFFFFFF0;
    // rom_array[40847] = 32'hFFFFFFF0;
    // rom_array[40848] = 32'hFFFFFFF0;
    // rom_array[40849] = 32'hFFFFFFF1;
    // rom_array[40850] = 32'hFFFFFFF1;
    // rom_array[40851] = 32'hFFFFFFF1;
    // rom_array[40852] = 32'hFFFFFFF1;
    // rom_array[40853] = 32'hFFFFFFF0;
    // rom_array[40854] = 32'hFFFFFFF0;
    // rom_array[40855] = 32'hFFFFFFF0;
    // rom_array[40856] = 32'hFFFFFFF0;
    // rom_array[40857] = 32'hFFFFFFF1;
    // rom_array[40858] = 32'hFFFFFFF1;
    // rom_array[40859] = 32'hFFFFFFF1;
    // rom_array[40860] = 32'hFFFFFFF1;
    // rom_array[40861] = 32'hFFFFFFF1;
    // rom_array[40862] = 32'hFFFFFFF1;
    // rom_array[40863] = 32'hFFFFFFF1;
    // rom_array[40864] = 32'hFFFFFFF1;
    // rom_array[40865] = 32'hFFFFFFF1;
    // rom_array[40866] = 32'hFFFFFFF1;
    // rom_array[40867] = 32'hFFFFFFF1;
    // rom_array[40868] = 32'hFFFFFFF1;
    // rom_array[40869] = 32'hFFFFFFF1;
    // rom_array[40870] = 32'hFFFFFFF1;
    // rom_array[40871] = 32'hFFFFFFF1;
    // rom_array[40872] = 32'hFFFFFFF1;
    // rom_array[40873] = 32'hFFFFFFF1;
    // rom_array[40874] = 32'hFFFFFFF1;
    // rom_array[40875] = 32'hFFFFFFF1;
    // rom_array[40876] = 32'hFFFFFFF1;
    // rom_array[40877] = 32'hFFFFFFF1;
    // rom_array[40878] = 32'hFFFFFFF1;
    // rom_array[40879] = 32'hFFFFFFF1;
    // rom_array[40880] = 32'hFFFFFFF1;
    // rom_array[40881] = 32'hFFFFFFF1;
    // rom_array[40882] = 32'hFFFFFFF1;
    // rom_array[40883] = 32'hFFFFFFF1;
    // rom_array[40884] = 32'hFFFFFFF1;
    // rom_array[40885] = 32'hFFFFFFF1;
    // rom_array[40886] = 32'hFFFFFFF1;
    // rom_array[40887] = 32'hFFFFFFF1;
    // rom_array[40888] = 32'hFFFFFFF1;
    // rom_array[40889] = 32'hFFFFFFF1;
    // rom_array[40890] = 32'hFFFFFFF1;
    // rom_array[40891] = 32'hFFFFFFF1;
    // rom_array[40892] = 32'hFFFFFFF1;
    // rom_array[40893] = 32'hFFFFFFF0;
    // rom_array[40894] = 32'hFFFFFFF0;
    // rom_array[40895] = 32'hFFFFFFF0;
    // rom_array[40896] = 32'hFFFFFFF0;
    // rom_array[40897] = 32'hFFFFFFF1;
    // rom_array[40898] = 32'hFFFFFFF1;
    // rom_array[40899] = 32'hFFFFFFF1;
    // rom_array[40900] = 32'hFFFFFFF1;
    // rom_array[40901] = 32'hFFFFFFF0;
    // rom_array[40902] = 32'hFFFFFFF0;
    // rom_array[40903] = 32'hFFFFFFF0;
    // rom_array[40904] = 32'hFFFFFFF0;
    // rom_array[40905] = 32'hFFFFFFF1;
    // rom_array[40906] = 32'hFFFFFFF1;
    // rom_array[40907] = 32'hFFFFFFF1;
    // rom_array[40908] = 32'hFFFFFFF1;
    // rom_array[40909] = 32'hFFFFFFF0;
    // rom_array[40910] = 32'hFFFFFFF0;
    // rom_array[40911] = 32'hFFFFFFF0;
    // rom_array[40912] = 32'hFFFFFFF0;
    // rom_array[40913] = 32'hFFFFFFF1;
    // rom_array[40914] = 32'hFFFFFFF1;
    // rom_array[40915] = 32'hFFFFFFF1;
    // rom_array[40916] = 32'hFFFFFFF1;
    // rom_array[40917] = 32'hFFFFFFF0;
    // rom_array[40918] = 32'hFFFFFFF0;
    // rom_array[40919] = 32'hFFFFFFF0;
    // rom_array[40920] = 32'hFFFFFFF0;
    // rom_array[40921] = 32'hFFFFFFF1;
    // rom_array[40922] = 32'hFFFFFFF1;
    // rom_array[40923] = 32'hFFFFFFF1;
    // rom_array[40924] = 32'hFFFFFFF1;
    // rom_array[40925] = 32'hFFFFFFF0;
    // rom_array[40926] = 32'hFFFFFFF0;
    // rom_array[40927] = 32'hFFFFFFF1;
    // rom_array[40928] = 32'hFFFFFFF1;
    // rom_array[40929] = 32'hFFFFFFF1;
    // rom_array[40930] = 32'hFFFFFFF1;
    // rom_array[40931] = 32'hFFFFFFF1;
    // rom_array[40932] = 32'hFFFFFFF1;
    // rom_array[40933] = 32'hFFFFFFF0;
    // rom_array[40934] = 32'hFFFFFFF0;
    // rom_array[40935] = 32'hFFFFFFF1;
    // rom_array[40936] = 32'hFFFFFFF1;
    // rom_array[40937] = 32'hFFFFFFF0;
    // rom_array[40938] = 32'hFFFFFFF0;
    // rom_array[40939] = 32'hFFFFFFF1;
    // rom_array[40940] = 32'hFFFFFFF1;
    // rom_array[40941] = 32'hFFFFFFF0;
    // rom_array[40942] = 32'hFFFFFFF0;
    // rom_array[40943] = 32'hFFFFFFF1;
    // rom_array[40944] = 32'hFFFFFFF1;
    // rom_array[40945] = 32'hFFFFFFF0;
    // rom_array[40946] = 32'hFFFFFFF0;
    // rom_array[40947] = 32'hFFFFFFF1;
    // rom_array[40948] = 32'hFFFFFFF1;
    // rom_array[40949] = 32'hFFFFFFF0;
    // rom_array[40950] = 32'hFFFFFFF0;
    // rom_array[40951] = 32'hFFFFFFF1;
    // rom_array[40952] = 32'hFFFFFFF1;
    // rom_array[40953] = 32'hFFFFFFF0;
    // rom_array[40954] = 32'hFFFFFFF0;
    // rom_array[40955] = 32'hFFFFFFF1;
    // rom_array[40956] = 32'hFFFFFFF1;
    // rom_array[40957] = 32'hFFFFFFF0;
    // rom_array[40958] = 32'hFFFFFFF0;
    // rom_array[40959] = 32'hFFFFFFF1;
    // rom_array[40960] = 32'hFFFFFFF1;
    // rom_array[40961] = 32'hFFFFFFF0;
    // rom_array[40962] = 32'hFFFFFFF0;
    // rom_array[40963] = 32'hFFFFFFF1;
    // rom_array[40964] = 32'hFFFFFFF1;
    // rom_array[40965] = 32'hFFFFFFF0;
    // rom_array[40966] = 32'hFFFFFFF0;
    // rom_array[40967] = 32'hFFFFFFF1;
    // rom_array[40968] = 32'hFFFFFFF1;
    // rom_array[40969] = 32'hFFFFFFF0;
    // rom_array[40970] = 32'hFFFFFFF0;
    // rom_array[40971] = 32'hFFFFFFF1;
    // rom_array[40972] = 32'hFFFFFFF1;
    // rom_array[40973] = 32'hFFFFFFF0;
    // rom_array[40974] = 32'hFFFFFFF0;
    // rom_array[40975] = 32'hFFFFFFF1;
    // rom_array[40976] = 32'hFFFFFFF1;
    // rom_array[40977] = 32'hFFFFFFF0;
    // rom_array[40978] = 32'hFFFFFFF0;
    // rom_array[40979] = 32'hFFFFFFF1;
    // rom_array[40980] = 32'hFFFFFFF1;
    // rom_array[40981] = 32'hFFFFFFF0;
    // rom_array[40982] = 32'hFFFFFFF0;
    // rom_array[40983] = 32'hFFFFFFF1;
    // rom_array[40984] = 32'hFFFFFFF1;
    // rom_array[40985] = 32'hFFFFFFF0;
    // rom_array[40986] = 32'hFFFFFFF0;
    // rom_array[40987] = 32'hFFFFFFF1;
    // rom_array[40988] = 32'hFFFFFFF1;
    // rom_array[40989] = 32'hFFFFFFF0;
    // rom_array[40990] = 32'hFFFFFFF0;
    // rom_array[40991] = 32'hFFFFFFF1;
    // rom_array[40992] = 32'hFFFFFFF1;
    // rom_array[40993] = 32'hFFFFFFF0;
    // rom_array[40994] = 32'hFFFFFFF0;
    // rom_array[40995] = 32'hFFFFFFF1;
    // rom_array[40996] = 32'hFFFFFFF1;
    // rom_array[40997] = 32'hFFFFFFF0;
    // rom_array[40998] = 32'hFFFFFFF0;
    // rom_array[40999] = 32'hFFFFFFF1;
    // rom_array[41000] = 32'hFFFFFFF1;
    // rom_array[41001] = 32'hFFFFFFF0;
    // rom_array[41002] = 32'hFFFFFFF0;
    // rom_array[41003] = 32'hFFFFFFF1;
    // rom_array[41004] = 32'hFFFFFFF1;
    // rom_array[41005] = 32'hFFFFFFF0;
    // rom_array[41006] = 32'hFFFFFFF0;
    // rom_array[41007] = 32'hFFFFFFF0;
    // rom_array[41008] = 32'hFFFFFFF0;
    // rom_array[41009] = 32'hFFFFFFF0;
    // rom_array[41010] = 32'hFFFFFFF0;
    // rom_array[41011] = 32'hFFFFFFF1;
    // rom_array[41012] = 32'hFFFFFFF1;
    // rom_array[41013] = 32'hFFFFFFF0;
    // rom_array[41014] = 32'hFFFFFFF0;
    // rom_array[41015] = 32'hFFFFFFF0;
    // rom_array[41016] = 32'hFFFFFFF0;
    // rom_array[41017] = 32'hFFFFFFF1;
    // rom_array[41018] = 32'hFFFFFFF1;
    // rom_array[41019] = 32'hFFFFFFF1;
    // rom_array[41020] = 32'hFFFFFFF1;
    // rom_array[41021] = 32'hFFFFFFF0;
    // rom_array[41022] = 32'hFFFFFFF0;
    // rom_array[41023] = 32'hFFFFFFF0;
    // rom_array[41024] = 32'hFFFFFFF0;
    // rom_array[41025] = 32'hFFFFFFF1;
    // rom_array[41026] = 32'hFFFFFFF1;
    // rom_array[41027] = 32'hFFFFFFF1;
    // rom_array[41028] = 32'hFFFFFFF1;
    // rom_array[41029] = 32'hFFFFFFF0;
    // rom_array[41030] = 32'hFFFFFFF0;
    // rom_array[41031] = 32'hFFFFFFF0;
    // rom_array[41032] = 32'hFFFFFFF0;
    // rom_array[41033] = 32'hFFFFFFF1;
    // rom_array[41034] = 32'hFFFFFFF1;
    // rom_array[41035] = 32'hFFFFFFF1;
    // rom_array[41036] = 32'hFFFFFFF1;
    // rom_array[41037] = 32'hFFFFFFF1;
    // rom_array[41038] = 32'hFFFFFFF1;
    // rom_array[41039] = 32'hFFFFFFF1;
    // rom_array[41040] = 32'hFFFFFFF1;
    // rom_array[41041] = 32'hFFFFFFF1;
    // rom_array[41042] = 32'hFFFFFFF1;
    // rom_array[41043] = 32'hFFFFFFF1;
    // rom_array[41044] = 32'hFFFFFFF1;
    // rom_array[41045] = 32'hFFFFFFF1;
    // rom_array[41046] = 32'hFFFFFFF1;
    // rom_array[41047] = 32'hFFFFFFF1;
    // rom_array[41048] = 32'hFFFFFFF1;
    // rom_array[41049] = 32'hFFFFFFF1;
    // rom_array[41050] = 32'hFFFFFFF1;
    // rom_array[41051] = 32'hFFFFFFF1;
    // rom_array[41052] = 32'hFFFFFFF1;
    // rom_array[41053] = 32'hFFFFFFF1;
    // rom_array[41054] = 32'hFFFFFFF1;
    // rom_array[41055] = 32'hFFFFFFF1;
    // rom_array[41056] = 32'hFFFFFFF1;
    // rom_array[41057] = 32'hFFFFFFF1;
    // rom_array[41058] = 32'hFFFFFFF1;
    // rom_array[41059] = 32'hFFFFFFF1;
    // rom_array[41060] = 32'hFFFFFFF1;
    // rom_array[41061] = 32'hFFFFFFF1;
    // rom_array[41062] = 32'hFFFFFFF1;
    // rom_array[41063] = 32'hFFFFFFF1;
    // rom_array[41064] = 32'hFFFFFFF1;
    // rom_array[41065] = 32'hFFFFFFF1;
    // rom_array[41066] = 32'hFFFFFFF1;
    // rom_array[41067] = 32'hFFFFFFF1;
    // rom_array[41068] = 32'hFFFFFFF1;
    // rom_array[41069] = 32'hFFFFFFF1;
    // rom_array[41070] = 32'hFFFFFFF1;
    // rom_array[41071] = 32'hFFFFFFF1;
    // rom_array[41072] = 32'hFFFFFFF1;
    // rom_array[41073] = 32'hFFFFFFF1;
    // rom_array[41074] = 32'hFFFFFFF1;
    // rom_array[41075] = 32'hFFFFFFF1;
    // rom_array[41076] = 32'hFFFFFFF1;
    // rom_array[41077] = 32'hFFFFFFF1;
    // rom_array[41078] = 32'hFFFFFFF1;
    // rom_array[41079] = 32'hFFFFFFF1;
    // rom_array[41080] = 32'hFFFFFFF1;
    // rom_array[41081] = 32'hFFFFFFF1;
    // rom_array[41082] = 32'hFFFFFFF1;
    // rom_array[41083] = 32'hFFFFFFF1;
    // rom_array[41084] = 32'hFFFFFFF1;
    // rom_array[41085] = 32'hFFFFFFF1;
    // rom_array[41086] = 32'hFFFFFFF1;
    // rom_array[41087] = 32'hFFFFFFF1;
    // rom_array[41088] = 32'hFFFFFFF1;
    // rom_array[41089] = 32'hFFFFFFF1;
    // rom_array[41090] = 32'hFFFFFFF1;
    // rom_array[41091] = 32'hFFFFFFF1;
    // rom_array[41092] = 32'hFFFFFFF1;
    // rom_array[41093] = 32'hFFFFFFF1;
    // rom_array[41094] = 32'hFFFFFFF1;
    // rom_array[41095] = 32'hFFFFFFF1;
    // rom_array[41096] = 32'hFFFFFFF1;
    // rom_array[41097] = 32'hFFFFFFF1;
    // rom_array[41098] = 32'hFFFFFFF1;
    // rom_array[41099] = 32'hFFFFFFF1;
    // rom_array[41100] = 32'hFFFFFFF1;
    // rom_array[41101] = 32'hFFFFFFF1;
    // rom_array[41102] = 32'hFFFFFFF1;
    // rom_array[41103] = 32'hFFFFFFF1;
    // rom_array[41104] = 32'hFFFFFFF1;
    // rom_array[41105] = 32'hFFFFFFF1;
    // rom_array[41106] = 32'hFFFFFFF1;
    // rom_array[41107] = 32'hFFFFFFF1;
    // rom_array[41108] = 32'hFFFFFFF1;
    // rom_array[41109] = 32'hFFFFFFF1;
    // rom_array[41110] = 32'hFFFFFFF1;
    // rom_array[41111] = 32'hFFFFFFF1;
    // rom_array[41112] = 32'hFFFFFFF1;
    // rom_array[41113] = 32'hFFFFFFF1;
    // rom_array[41114] = 32'hFFFFFFF1;
    // rom_array[41115] = 32'hFFFFFFF1;
    // rom_array[41116] = 32'hFFFFFFF1;
    // rom_array[41117] = 32'hFFFFFFF1;
    // rom_array[41118] = 32'hFFFFFFF1;
    // rom_array[41119] = 32'hFFFFFFF1;
    // rom_array[41120] = 32'hFFFFFFF1;
    // rom_array[41121] = 32'hFFFFFFF1;
    // rom_array[41122] = 32'hFFFFFFF1;
    // rom_array[41123] = 32'hFFFFFFF1;
    // rom_array[41124] = 32'hFFFFFFF1;
    // rom_array[41125] = 32'hFFFFFFF1;
    // rom_array[41126] = 32'hFFFFFFF1;
    // rom_array[41127] = 32'hFFFFFFF1;
    // rom_array[41128] = 32'hFFFFFFF1;
    // rom_array[41129] = 32'hFFFFFFF1;
    // rom_array[41130] = 32'hFFFFFFF1;
    // rom_array[41131] = 32'hFFFFFFF1;
    // rom_array[41132] = 32'hFFFFFFF1;
    // rom_array[41133] = 32'hFFFFFFF0;
    // rom_array[41134] = 32'hFFFFFFF0;
    // rom_array[41135] = 32'hFFFFFFF0;
    // rom_array[41136] = 32'hFFFFFFF0;
    // rom_array[41137] = 32'hFFFFFFF1;
    // rom_array[41138] = 32'hFFFFFFF1;
    // rom_array[41139] = 32'hFFFFFFF1;
    // rom_array[41140] = 32'hFFFFFFF1;
    // rom_array[41141] = 32'hFFFFFFF0;
    // rom_array[41142] = 32'hFFFFFFF0;
    // rom_array[41143] = 32'hFFFFFFF0;
    // rom_array[41144] = 32'hFFFFFFF0;
    // rom_array[41145] = 32'hFFFFFFF1;
    // rom_array[41146] = 32'hFFFFFFF1;
    // rom_array[41147] = 32'hFFFFFFF1;
    // rom_array[41148] = 32'hFFFFFFF1;
    // rom_array[41149] = 32'hFFFFFFF0;
    // rom_array[41150] = 32'hFFFFFFF0;
    // rom_array[41151] = 32'hFFFFFFF0;
    // rom_array[41152] = 32'hFFFFFFF0;
    // rom_array[41153] = 32'hFFFFFFF1;
    // rom_array[41154] = 32'hFFFFFFF1;
    // rom_array[41155] = 32'hFFFFFFF1;
    // rom_array[41156] = 32'hFFFFFFF1;
    // rom_array[41157] = 32'hFFFFFFF0;
    // rom_array[41158] = 32'hFFFFFFF0;
    // rom_array[41159] = 32'hFFFFFFF0;
    // rom_array[41160] = 32'hFFFFFFF0;
    // rom_array[41161] = 32'hFFFFFFF1;
    // rom_array[41162] = 32'hFFFFFFF1;
    // rom_array[41163] = 32'hFFFFFFF1;
    // rom_array[41164] = 32'hFFFFFFF1;
    // rom_array[41165] = 32'hFFFFFFF1;
    // rom_array[41166] = 32'hFFFFFFF1;
    // rom_array[41167] = 32'hFFFFFFF1;
    // rom_array[41168] = 32'hFFFFFFF1;
    // rom_array[41169] = 32'hFFFFFFF1;
    // rom_array[41170] = 32'hFFFFFFF1;
    // rom_array[41171] = 32'hFFFFFFF1;
    // rom_array[41172] = 32'hFFFFFFF1;
    // rom_array[41173] = 32'hFFFFFFF1;
    // rom_array[41174] = 32'hFFFFFFF1;
    // rom_array[41175] = 32'hFFFFFFF1;
    // rom_array[41176] = 32'hFFFFFFF1;
    // rom_array[41177] = 32'hFFFFFFF1;
    // rom_array[41178] = 32'hFFFFFFF1;
    // rom_array[41179] = 32'hFFFFFFF1;
    // rom_array[41180] = 32'hFFFFFFF1;
    // rom_array[41181] = 32'hFFFFFFF0;
    // rom_array[41182] = 32'hFFFFFFF0;
    // rom_array[41183] = 32'hFFFFFFF0;
    // rom_array[41184] = 32'hFFFFFFF0;
    // rom_array[41185] = 32'hFFFFFFF1;
    // rom_array[41186] = 32'hFFFFFFF1;
    // rom_array[41187] = 32'hFFFFFFF1;
    // rom_array[41188] = 32'hFFFFFFF1;
    // rom_array[41189] = 32'hFFFFFFF0;
    // rom_array[41190] = 32'hFFFFFFF0;
    // rom_array[41191] = 32'hFFFFFFF0;
    // rom_array[41192] = 32'hFFFFFFF0;
    // rom_array[41193] = 32'hFFFFFFF0;
    // rom_array[41194] = 32'hFFFFFFF0;
    // rom_array[41195] = 32'hFFFFFFF0;
    // rom_array[41196] = 32'hFFFFFFF0;
    // rom_array[41197] = 32'hFFFFFFF1;
    // rom_array[41198] = 32'hFFFFFFF1;
    // rom_array[41199] = 32'hFFFFFFF1;
    // rom_array[41200] = 32'hFFFFFFF1;
    // rom_array[41201] = 32'hFFFFFFF0;
    // rom_array[41202] = 32'hFFFFFFF0;
    // rom_array[41203] = 32'hFFFFFFF0;
    // rom_array[41204] = 32'hFFFFFFF0;
    // rom_array[41205] = 32'hFFFFFFF1;
    // rom_array[41206] = 32'hFFFFFFF1;
    // rom_array[41207] = 32'hFFFFFFF1;
    // rom_array[41208] = 32'hFFFFFFF1;
    // rom_array[41209] = 32'hFFFFFFF0;
    // rom_array[41210] = 32'hFFFFFFF0;
    // rom_array[41211] = 32'hFFFFFFF0;
    // rom_array[41212] = 32'hFFFFFFF0;
    // rom_array[41213] = 32'hFFFFFFF1;
    // rom_array[41214] = 32'hFFFFFFF1;
    // rom_array[41215] = 32'hFFFFFFF1;
    // rom_array[41216] = 32'hFFFFFFF1;
    // rom_array[41217] = 32'hFFFFFFF0;
    // rom_array[41218] = 32'hFFFFFFF0;
    // rom_array[41219] = 32'hFFFFFFF0;
    // rom_array[41220] = 32'hFFFFFFF0;
    // rom_array[41221] = 32'hFFFFFFF1;
    // rom_array[41222] = 32'hFFFFFFF1;
    // rom_array[41223] = 32'hFFFFFFF1;
    // rom_array[41224] = 32'hFFFFFFF1;
    // rom_array[41225] = 32'hFFFFFFF0;
    // rom_array[41226] = 32'hFFFFFFF0;
    // rom_array[41227] = 32'hFFFFFFF0;
    // rom_array[41228] = 32'hFFFFFFF0;
    // rom_array[41229] = 32'hFFFFFFF1;
    // rom_array[41230] = 32'hFFFFFFF1;
    // rom_array[41231] = 32'hFFFFFFF1;
    // rom_array[41232] = 32'hFFFFFFF1;
    // rom_array[41233] = 32'hFFFFFFF0;
    // rom_array[41234] = 32'hFFFFFFF0;
    // rom_array[41235] = 32'hFFFFFFF0;
    // rom_array[41236] = 32'hFFFFFFF0;
    // rom_array[41237] = 32'hFFFFFFF1;
    // rom_array[41238] = 32'hFFFFFFF1;
    // rom_array[41239] = 32'hFFFFFFF1;
    // rom_array[41240] = 32'hFFFFFFF1;
    // rom_array[41241] = 32'hFFFFFFF0;
    // rom_array[41242] = 32'hFFFFFFF0;
    // rom_array[41243] = 32'hFFFFFFF0;
    // rom_array[41244] = 32'hFFFFFFF0;
    // rom_array[41245] = 32'hFFFFFFF1;
    // rom_array[41246] = 32'hFFFFFFF1;
    // rom_array[41247] = 32'hFFFFFFF1;
    // rom_array[41248] = 32'hFFFFFFF1;
    // rom_array[41249] = 32'hFFFFFFF0;
    // rom_array[41250] = 32'hFFFFFFF0;
    // rom_array[41251] = 32'hFFFFFFF0;
    // rom_array[41252] = 32'hFFFFFFF0;
    // rom_array[41253] = 32'hFFFFFFF1;
    // rom_array[41254] = 32'hFFFFFFF1;
    // rom_array[41255] = 32'hFFFFFFF1;
    // rom_array[41256] = 32'hFFFFFFF1;
    // rom_array[41257] = 32'hFFFFFFF0;
    // rom_array[41258] = 32'hFFFFFFF0;
    // rom_array[41259] = 32'hFFFFFFF0;
    // rom_array[41260] = 32'hFFFFFFF0;
    // rom_array[41261] = 32'hFFFFFFF1;
    // rom_array[41262] = 32'hFFFFFFF1;
    // rom_array[41263] = 32'hFFFFFFF1;
    // rom_array[41264] = 32'hFFFFFFF1;
    // rom_array[41265] = 32'hFFFFFFF0;
    // rom_array[41266] = 32'hFFFFFFF0;
    // rom_array[41267] = 32'hFFFFFFF0;
    // rom_array[41268] = 32'hFFFFFFF0;
    // rom_array[41269] = 32'hFFFFFFF1;
    // rom_array[41270] = 32'hFFFFFFF1;
    // rom_array[41271] = 32'hFFFFFFF1;
    // rom_array[41272] = 32'hFFFFFFF1;
    // rom_array[41273] = 32'hFFFFFFF0;
    // rom_array[41274] = 32'hFFFFFFF0;
    // rom_array[41275] = 32'hFFFFFFF0;
    // rom_array[41276] = 32'hFFFFFFF0;
    // rom_array[41277] = 32'hFFFFFFF1;
    // rom_array[41278] = 32'hFFFFFFF1;
    // rom_array[41279] = 32'hFFFFFFF1;
    // rom_array[41280] = 32'hFFFFFFF1;
    // rom_array[41281] = 32'hFFFFFFF0;
    // rom_array[41282] = 32'hFFFFFFF0;
    // rom_array[41283] = 32'hFFFFFFF0;
    // rom_array[41284] = 32'hFFFFFFF0;
    // rom_array[41285] = 32'hFFFFFFF1;
    // rom_array[41286] = 32'hFFFFFFF1;
    // rom_array[41287] = 32'hFFFFFFF1;
    // rom_array[41288] = 32'hFFFFFFF1;
    // rom_array[41289] = 32'hFFFFFFF0;
    // rom_array[41290] = 32'hFFFFFFF0;
    // rom_array[41291] = 32'hFFFFFFF0;
    // rom_array[41292] = 32'hFFFFFFF0;
    // rom_array[41293] = 32'hFFFFFFF1;
    // rom_array[41294] = 32'hFFFFFFF1;
    // rom_array[41295] = 32'hFFFFFFF1;
    // rom_array[41296] = 32'hFFFFFFF1;
    // rom_array[41297] = 32'hFFFFFFF0;
    // rom_array[41298] = 32'hFFFFFFF0;
    // rom_array[41299] = 32'hFFFFFFF0;
    // rom_array[41300] = 32'hFFFFFFF0;
    // rom_array[41301] = 32'hFFFFFFF1;
    // rom_array[41302] = 32'hFFFFFFF1;
    // rom_array[41303] = 32'hFFFFFFF1;
    // rom_array[41304] = 32'hFFFFFFF1;
    // rom_array[41305] = 32'hFFFFFFF0;
    // rom_array[41306] = 32'hFFFFFFF0;
    // rom_array[41307] = 32'hFFFFFFF0;
    // rom_array[41308] = 32'hFFFFFFF0;
    // rom_array[41309] = 32'hFFFFFFF1;
    // rom_array[41310] = 32'hFFFFFFF1;
    // rom_array[41311] = 32'hFFFFFFF1;
    // rom_array[41312] = 32'hFFFFFFF1;
    // rom_array[41313] = 32'hFFFFFFF0;
    // rom_array[41314] = 32'hFFFFFFF0;
    // rom_array[41315] = 32'hFFFFFFF0;
    // rom_array[41316] = 32'hFFFFFFF0;
    // rom_array[41317] = 32'hFFFFFFF1;
    // rom_array[41318] = 32'hFFFFFFF1;
    // rom_array[41319] = 32'hFFFFFFF1;
    // rom_array[41320] = 32'hFFFFFFF1;
    // rom_array[41321] = 32'hFFFFFFF0;
    // rom_array[41322] = 32'hFFFFFFF0;
    // rom_array[41323] = 32'hFFFFFFF0;
    // rom_array[41324] = 32'hFFFFFFF0;
    // rom_array[41325] = 32'hFFFFFFF1;
    // rom_array[41326] = 32'hFFFFFFF1;
    // rom_array[41327] = 32'hFFFFFFF1;
    // rom_array[41328] = 32'hFFFFFFF1;
    // rom_array[41329] = 32'hFFFFFFF0;
    // rom_array[41330] = 32'hFFFFFFF0;
    // rom_array[41331] = 32'hFFFFFFF0;
    // rom_array[41332] = 32'hFFFFFFF0;
    // rom_array[41333] = 32'hFFFFFFF1;
    // rom_array[41334] = 32'hFFFFFFF1;
    // rom_array[41335] = 32'hFFFFFFF1;
    // rom_array[41336] = 32'hFFFFFFF1;
    // rom_array[41337] = 32'hFFFFFFF0;
    // rom_array[41338] = 32'hFFFFFFF0;
    // rom_array[41339] = 32'hFFFFFFF0;
    // rom_array[41340] = 32'hFFFFFFF0;
    // rom_array[41341] = 32'hFFFFFFF1;
    // rom_array[41342] = 32'hFFFFFFF1;
    // rom_array[41343] = 32'hFFFFFFF1;
    // rom_array[41344] = 32'hFFFFFFF1;
    // rom_array[41345] = 32'hFFFFFFF0;
    // rom_array[41346] = 32'hFFFFFFF0;
    // rom_array[41347] = 32'hFFFFFFF0;
    // rom_array[41348] = 32'hFFFFFFF0;
    // rom_array[41349] = 32'hFFFFFFF1;
    // rom_array[41350] = 32'hFFFFFFF1;
    // rom_array[41351] = 32'hFFFFFFF1;
    // rom_array[41352] = 32'hFFFFFFF1;
    // rom_array[41353] = 32'hFFFFFFF0;
    // rom_array[41354] = 32'hFFFFFFF0;
    // rom_array[41355] = 32'hFFFFFFF0;
    // rom_array[41356] = 32'hFFFFFFF0;
    // rom_array[41357] = 32'hFFFFFFF1;
    // rom_array[41358] = 32'hFFFFFFF1;
    // rom_array[41359] = 32'hFFFFFFF1;
    // rom_array[41360] = 32'hFFFFFFF1;
    // rom_array[41361] = 32'hFFFFFFF0;
    // rom_array[41362] = 32'hFFFFFFF0;
    // rom_array[41363] = 32'hFFFFFFF0;
    // rom_array[41364] = 32'hFFFFFFF0;
    // rom_array[41365] = 32'hFFFFFFF1;
    // rom_array[41366] = 32'hFFFFFFF1;
    // rom_array[41367] = 32'hFFFFFFF1;
    // rom_array[41368] = 32'hFFFFFFF1;
    // rom_array[41369] = 32'hFFFFFFF1;
    // rom_array[41370] = 32'hFFFFFFF1;
    // rom_array[41371] = 32'hFFFFFFF1;
    // rom_array[41372] = 32'hFFFFFFF1;
    // rom_array[41373] = 32'hFFFFFFF1;
    // rom_array[41374] = 32'hFFFFFFF1;
    // rom_array[41375] = 32'hFFFFFFF1;
    // rom_array[41376] = 32'hFFFFFFF1;
    // rom_array[41377] = 32'hFFFFFFF1;
    // rom_array[41378] = 32'hFFFFFFF1;
    // rom_array[41379] = 32'hFFFFFFF1;
    // rom_array[41380] = 32'hFFFFFFF1;
    // rom_array[41381] = 32'hFFFFFFF1;
    // rom_array[41382] = 32'hFFFFFFF1;
    // rom_array[41383] = 32'hFFFFFFF1;
    // rom_array[41384] = 32'hFFFFFFF1;
    // rom_array[41385] = 32'hFFFFFFF1;
    // rom_array[41386] = 32'hFFFFFFF1;
    // rom_array[41387] = 32'hFFFFFFF1;
    // rom_array[41388] = 32'hFFFFFFF1;
    // rom_array[41389] = 32'hFFFFFFF1;
    // rom_array[41390] = 32'hFFFFFFF1;
    // rom_array[41391] = 32'hFFFFFFF1;
    // rom_array[41392] = 32'hFFFFFFF1;
    // rom_array[41393] = 32'hFFFFFFF1;
    // rom_array[41394] = 32'hFFFFFFF1;
    // rom_array[41395] = 32'hFFFFFFF1;
    // rom_array[41396] = 32'hFFFFFFF1;
    // rom_array[41397] = 32'hFFFFFFF1;
    // rom_array[41398] = 32'hFFFFFFF1;
    // rom_array[41399] = 32'hFFFFFFF1;
    // rom_array[41400] = 32'hFFFFFFF1;
    // rom_array[41401] = 32'hFFFFFFF1;
    // rom_array[41402] = 32'hFFFFFFF1;
    // rom_array[41403] = 32'hFFFFFFF1;
    // rom_array[41404] = 32'hFFFFFFF1;
    // rom_array[41405] = 32'hFFFFFFF1;
    // rom_array[41406] = 32'hFFFFFFF1;
    // rom_array[41407] = 32'hFFFFFFF1;
    // rom_array[41408] = 32'hFFFFFFF1;
    // rom_array[41409] = 32'hFFFFFFF1;
    // rom_array[41410] = 32'hFFFFFFF1;
    // rom_array[41411] = 32'hFFFFFFF1;
    // rom_array[41412] = 32'hFFFFFFF1;
    // rom_array[41413] = 32'hFFFFFFF1;
    // rom_array[41414] = 32'hFFFFFFF1;
    // rom_array[41415] = 32'hFFFFFFF1;
    // rom_array[41416] = 32'hFFFFFFF1;
    // rom_array[41417] = 32'hFFFFFFF1;
    // rom_array[41418] = 32'hFFFFFFF1;
    // rom_array[41419] = 32'hFFFFFFF1;
    // rom_array[41420] = 32'hFFFFFFF1;
    // rom_array[41421] = 32'hFFFFFFF1;
    // rom_array[41422] = 32'hFFFFFFF1;
    // rom_array[41423] = 32'hFFFFFFF1;
    // rom_array[41424] = 32'hFFFFFFF1;
    // rom_array[41425] = 32'hFFFFFFF1;
    // rom_array[41426] = 32'hFFFFFFF1;
    // rom_array[41427] = 32'hFFFFFFF1;
    // rom_array[41428] = 32'hFFFFFFF1;
    // rom_array[41429] = 32'hFFFFFFF1;
    // rom_array[41430] = 32'hFFFFFFF1;
    // rom_array[41431] = 32'hFFFFFFF1;
    // rom_array[41432] = 32'hFFFFFFF1;
    // rom_array[41433] = 32'hFFFFFFF1;
    // rom_array[41434] = 32'hFFFFFFF1;
    // rom_array[41435] = 32'hFFFFFFF1;
    // rom_array[41436] = 32'hFFFFFFF1;
    // rom_array[41437] = 32'hFFFFFFF1;
    // rom_array[41438] = 32'hFFFFFFF1;
    // rom_array[41439] = 32'hFFFFFFF1;
    // rom_array[41440] = 32'hFFFFFFF1;
    // rom_array[41441] = 32'hFFFFFFF1;
    // rom_array[41442] = 32'hFFFFFFF1;
    // rom_array[41443] = 32'hFFFFFFF1;
    // rom_array[41444] = 32'hFFFFFFF1;
    // rom_array[41445] = 32'hFFFFFFF1;
    // rom_array[41446] = 32'hFFFFFFF1;
    // rom_array[41447] = 32'hFFFFFFF1;
    // rom_array[41448] = 32'hFFFFFFF1;
    // rom_array[41449] = 32'hFFFFFFF1;
    // rom_array[41450] = 32'hFFFFFFF1;
    // rom_array[41451] = 32'hFFFFFFF1;
    // rom_array[41452] = 32'hFFFFFFF1;
    // rom_array[41453] = 32'hFFFFFFF1;
    // rom_array[41454] = 32'hFFFFFFF1;
    // rom_array[41455] = 32'hFFFFFFF1;
    // rom_array[41456] = 32'hFFFFFFF1;
    // rom_array[41457] = 32'hFFFFFFF1;
    // rom_array[41458] = 32'hFFFFFFF1;
    // rom_array[41459] = 32'hFFFFFFF1;
    // rom_array[41460] = 32'hFFFFFFF1;
    // rom_array[41461] = 32'hFFFFFFF1;
    // rom_array[41462] = 32'hFFFFFFF1;
    // rom_array[41463] = 32'hFFFFFFF1;
    // rom_array[41464] = 32'hFFFFFFF1;
    // rom_array[41465] = 32'hFFFFFFF1;
    // rom_array[41466] = 32'hFFFFFFF1;
    // rom_array[41467] = 32'hFFFFFFF1;
    // rom_array[41468] = 32'hFFFFFFF1;
    // rom_array[41469] = 32'hFFFFFFF1;
    // rom_array[41470] = 32'hFFFFFFF1;
    // rom_array[41471] = 32'hFFFFFFF1;
    // rom_array[41472] = 32'hFFFFFFF1;
    // rom_array[41473] = 32'hFFFFFFF1;
    // rom_array[41474] = 32'hFFFFFFF1;
    // rom_array[41475] = 32'hFFFFFFF1;
    // rom_array[41476] = 32'hFFFFFFF1;
    // rom_array[41477] = 32'hFFFFFFF1;
    // rom_array[41478] = 32'hFFFFFFF1;
    // rom_array[41479] = 32'hFFFFFFF1;
    // rom_array[41480] = 32'hFFFFFFF1;
    // rom_array[41481] = 32'hFFFFFFF0;
    // rom_array[41482] = 32'hFFFFFFF0;
    // rom_array[41483] = 32'hFFFFFFF0;
    // rom_array[41484] = 32'hFFFFFFF0;
    // rom_array[41485] = 32'hFFFFFFF1;
    // rom_array[41486] = 32'hFFFFFFF1;
    // rom_array[41487] = 32'hFFFFFFF1;
    // rom_array[41488] = 32'hFFFFFFF1;
    // rom_array[41489] = 32'hFFFFFFF0;
    // rom_array[41490] = 32'hFFFFFFF0;
    // rom_array[41491] = 32'hFFFFFFF0;
    // rom_array[41492] = 32'hFFFFFFF0;
    // rom_array[41493] = 32'hFFFFFFF1;
    // rom_array[41494] = 32'hFFFFFFF1;
    // rom_array[41495] = 32'hFFFFFFF1;
    // rom_array[41496] = 32'hFFFFFFF1;
    // rom_array[41497] = 32'hFFFFFFF0;
    // rom_array[41498] = 32'hFFFFFFF0;
    // rom_array[41499] = 32'hFFFFFFF0;
    // rom_array[41500] = 32'hFFFFFFF0;
    // rom_array[41501] = 32'hFFFFFFF1;
    // rom_array[41502] = 32'hFFFFFFF1;
    // rom_array[41503] = 32'hFFFFFFF1;
    // rom_array[41504] = 32'hFFFFFFF1;
    // rom_array[41505] = 32'hFFFFFFF0;
    // rom_array[41506] = 32'hFFFFFFF0;
    // rom_array[41507] = 32'hFFFFFFF0;
    // rom_array[41508] = 32'hFFFFFFF0;
    // rom_array[41509] = 32'hFFFFFFF1;
    // rom_array[41510] = 32'hFFFFFFF1;
    // rom_array[41511] = 32'hFFFFFFF1;
    // rom_array[41512] = 32'hFFFFFFF1;
    // rom_array[41513] = 32'hFFFFFFF0;
    // rom_array[41514] = 32'hFFFFFFF0;
    // rom_array[41515] = 32'hFFFFFFF0;
    // rom_array[41516] = 32'hFFFFFFF0;
    // rom_array[41517] = 32'hFFFFFFF1;
    // rom_array[41518] = 32'hFFFFFFF1;
    // rom_array[41519] = 32'hFFFFFFF1;
    // rom_array[41520] = 32'hFFFFFFF1;
    // rom_array[41521] = 32'hFFFFFFF0;
    // rom_array[41522] = 32'hFFFFFFF0;
    // rom_array[41523] = 32'hFFFFFFF0;
    // rom_array[41524] = 32'hFFFFFFF0;
    // rom_array[41525] = 32'hFFFFFFF1;
    // rom_array[41526] = 32'hFFFFFFF1;
    // rom_array[41527] = 32'hFFFFFFF1;
    // rom_array[41528] = 32'hFFFFFFF1;
    // rom_array[41529] = 32'hFFFFFFF0;
    // rom_array[41530] = 32'hFFFFFFF0;
    // rom_array[41531] = 32'hFFFFFFF0;
    // rom_array[41532] = 32'hFFFFFFF0;
    // rom_array[41533] = 32'hFFFFFFF1;
    // rom_array[41534] = 32'hFFFFFFF1;
    // rom_array[41535] = 32'hFFFFFFF1;
    // rom_array[41536] = 32'hFFFFFFF1;
    // rom_array[41537] = 32'hFFFFFFF0;
    // rom_array[41538] = 32'hFFFFFFF0;
    // rom_array[41539] = 32'hFFFFFFF0;
    // rom_array[41540] = 32'hFFFFFFF0;
    // rom_array[41541] = 32'hFFFFFFF1;
    // rom_array[41542] = 32'hFFFFFFF1;
    // rom_array[41543] = 32'hFFFFFFF1;
    // rom_array[41544] = 32'hFFFFFFF1;
    // rom_array[41545] = 32'hFFFFFFF0;
    // rom_array[41546] = 32'hFFFFFFF0;
    // rom_array[41547] = 32'hFFFFFFF0;
    // rom_array[41548] = 32'hFFFFFFF0;
    // rom_array[41549] = 32'hFFFFFFF1;
    // rom_array[41550] = 32'hFFFFFFF1;
    // rom_array[41551] = 32'hFFFFFFF1;
    // rom_array[41552] = 32'hFFFFFFF1;
    // rom_array[41553] = 32'hFFFFFFF0;
    // rom_array[41554] = 32'hFFFFFFF0;
    // rom_array[41555] = 32'hFFFFFFF0;
    // rom_array[41556] = 32'hFFFFFFF0;
    // rom_array[41557] = 32'hFFFFFFF1;
    // rom_array[41558] = 32'hFFFFFFF1;
    // rom_array[41559] = 32'hFFFFFFF1;
    // rom_array[41560] = 32'hFFFFFFF1;
    // rom_array[41561] = 32'hFFFFFFF0;
    // rom_array[41562] = 32'hFFFFFFF0;
    // rom_array[41563] = 32'hFFFFFFF0;
    // rom_array[41564] = 32'hFFFFFFF0;
    // rom_array[41565] = 32'hFFFFFFF1;
    // rom_array[41566] = 32'hFFFFFFF1;
    // rom_array[41567] = 32'hFFFFFFF1;
    // rom_array[41568] = 32'hFFFFFFF1;
    // rom_array[41569] = 32'hFFFFFFF0;
    // rom_array[41570] = 32'hFFFFFFF0;
    // rom_array[41571] = 32'hFFFFFFF0;
    // rom_array[41572] = 32'hFFFFFFF0;
    // rom_array[41573] = 32'hFFFFFFF1;
    // rom_array[41574] = 32'hFFFFFFF1;
    // rom_array[41575] = 32'hFFFFFFF1;
    // rom_array[41576] = 32'hFFFFFFF1;
    // rom_array[41577] = 32'hFFFFFFF0;
    // rom_array[41578] = 32'hFFFFFFF0;
    // rom_array[41579] = 32'hFFFFFFF0;
    // rom_array[41580] = 32'hFFFFFFF0;
    // rom_array[41581] = 32'hFFFFFFF1;
    // rom_array[41582] = 32'hFFFFFFF1;
    // rom_array[41583] = 32'hFFFFFFF1;
    // rom_array[41584] = 32'hFFFFFFF1;
    // rom_array[41585] = 32'hFFFFFFF0;
    // rom_array[41586] = 32'hFFFFFFF0;
    // rom_array[41587] = 32'hFFFFFFF0;
    // rom_array[41588] = 32'hFFFFFFF0;
    // rom_array[41589] = 32'hFFFFFFF1;
    // rom_array[41590] = 32'hFFFFFFF1;
    // rom_array[41591] = 32'hFFFFFFF1;
    // rom_array[41592] = 32'hFFFFFFF1;
    // rom_array[41593] = 32'hFFFFFFF0;
    // rom_array[41594] = 32'hFFFFFFF0;
    // rom_array[41595] = 32'hFFFFFFF0;
    // rom_array[41596] = 32'hFFFFFFF0;
    // rom_array[41597] = 32'hFFFFFFF1;
    // rom_array[41598] = 32'hFFFFFFF1;
    // rom_array[41599] = 32'hFFFFFFF1;
    // rom_array[41600] = 32'hFFFFFFF1;
    // rom_array[41601] = 32'hFFFFFFF0;
    // rom_array[41602] = 32'hFFFFFFF0;
    // rom_array[41603] = 32'hFFFFFFF0;
    // rom_array[41604] = 32'hFFFFFFF0;
    // rom_array[41605] = 32'hFFFFFFF1;
    // rom_array[41606] = 32'hFFFFFFF1;
    // rom_array[41607] = 32'hFFFFFFF1;
    // rom_array[41608] = 32'hFFFFFFF1;
    // rom_array[41609] = 32'hFFFFFFF0;
    // rom_array[41610] = 32'hFFFFFFF0;
    // rom_array[41611] = 32'hFFFFFFF1;
    // rom_array[41612] = 32'hFFFFFFF1;
    // rom_array[41613] = 32'hFFFFFFF0;
    // rom_array[41614] = 32'hFFFFFFF0;
    // rom_array[41615] = 32'hFFFFFFF1;
    // rom_array[41616] = 32'hFFFFFFF1;
    // rom_array[41617] = 32'hFFFFFFF0;
    // rom_array[41618] = 32'hFFFFFFF0;
    // rom_array[41619] = 32'hFFFFFFF1;
    // rom_array[41620] = 32'hFFFFFFF1;
    // rom_array[41621] = 32'hFFFFFFF0;
    // rom_array[41622] = 32'hFFFFFFF0;
    // rom_array[41623] = 32'hFFFFFFF1;
    // rom_array[41624] = 32'hFFFFFFF1;
    // rom_array[41625] = 32'hFFFFFFF0;
    // rom_array[41626] = 32'hFFFFFFF0;
    // rom_array[41627] = 32'hFFFFFFF1;
    // rom_array[41628] = 32'hFFFFFFF1;
    // rom_array[41629] = 32'hFFFFFFF0;
    // rom_array[41630] = 32'hFFFFFFF0;
    // rom_array[41631] = 32'hFFFFFFF1;
    // rom_array[41632] = 32'hFFFFFFF1;
    // rom_array[41633] = 32'hFFFFFFF0;
    // rom_array[41634] = 32'hFFFFFFF0;
    // rom_array[41635] = 32'hFFFFFFF1;
    // rom_array[41636] = 32'hFFFFFFF1;
    // rom_array[41637] = 32'hFFFFFFF0;
    // rom_array[41638] = 32'hFFFFFFF0;
    // rom_array[41639] = 32'hFFFFFFF1;
    // rom_array[41640] = 32'hFFFFFFF1;
    // rom_array[41641] = 32'hFFFFFFF0;
    // rom_array[41642] = 32'hFFFFFFF0;
    // rom_array[41643] = 32'hFFFFFFF1;
    // rom_array[41644] = 32'hFFFFFFF1;
    // rom_array[41645] = 32'hFFFFFFF0;
    // rom_array[41646] = 32'hFFFFFFF0;
    // rom_array[41647] = 32'hFFFFFFF1;
    // rom_array[41648] = 32'hFFFFFFF1;
    // rom_array[41649] = 32'hFFFFFFF0;
    // rom_array[41650] = 32'hFFFFFFF0;
    // rom_array[41651] = 32'hFFFFFFF1;
    // rom_array[41652] = 32'hFFFFFFF1;
    // rom_array[41653] = 32'hFFFFFFF0;
    // rom_array[41654] = 32'hFFFFFFF0;
    // rom_array[41655] = 32'hFFFFFFF1;
    // rom_array[41656] = 32'hFFFFFFF1;
    // rom_array[41657] = 32'hFFFFFFF1;
    // rom_array[41658] = 32'hFFFFFFF1;
    // rom_array[41659] = 32'hFFFFFFF1;
    // rom_array[41660] = 32'hFFFFFFF1;
    // rom_array[41661] = 32'hFFFFFFF0;
    // rom_array[41662] = 32'hFFFFFFF0;
    // rom_array[41663] = 32'hFFFFFFF0;
    // rom_array[41664] = 32'hFFFFFFF0;
    // rom_array[41665] = 32'hFFFFFFF1;
    // rom_array[41666] = 32'hFFFFFFF1;
    // rom_array[41667] = 32'hFFFFFFF1;
    // rom_array[41668] = 32'hFFFFFFF1;
    // rom_array[41669] = 32'hFFFFFFF0;
    // rom_array[41670] = 32'hFFFFFFF0;
    // rom_array[41671] = 32'hFFFFFFF0;
    // rom_array[41672] = 32'hFFFFFFF0;
    // rom_array[41673] = 32'hFFFFFFF1;
    // rom_array[41674] = 32'hFFFFFFF1;
    // rom_array[41675] = 32'hFFFFFFF1;
    // rom_array[41676] = 32'hFFFFFFF1;
    // rom_array[41677] = 32'hFFFFFFF0;
    // rom_array[41678] = 32'hFFFFFFF0;
    // rom_array[41679] = 32'hFFFFFFF0;
    // rom_array[41680] = 32'hFFFFFFF0;
    // rom_array[41681] = 32'hFFFFFFF1;
    // rom_array[41682] = 32'hFFFFFFF1;
    // rom_array[41683] = 32'hFFFFFFF1;
    // rom_array[41684] = 32'hFFFFFFF1;
    // rom_array[41685] = 32'hFFFFFFF0;
    // rom_array[41686] = 32'hFFFFFFF0;
    // rom_array[41687] = 32'hFFFFFFF0;
    // rom_array[41688] = 32'hFFFFFFF0;
    // rom_array[41689] = 32'hFFFFFFF1;
    // rom_array[41690] = 32'hFFFFFFF1;
    // rom_array[41691] = 32'hFFFFFFF1;
    // rom_array[41692] = 32'hFFFFFFF1;
    // rom_array[41693] = 32'hFFFFFFF0;
    // rom_array[41694] = 32'hFFFFFFF0;
    // rom_array[41695] = 32'hFFFFFFF0;
    // rom_array[41696] = 32'hFFFFFFF0;
    // rom_array[41697] = 32'hFFFFFFF1;
    // rom_array[41698] = 32'hFFFFFFF1;
    // rom_array[41699] = 32'hFFFFFFF1;
    // rom_array[41700] = 32'hFFFFFFF1;
    // rom_array[41701] = 32'hFFFFFFF0;
    // rom_array[41702] = 32'hFFFFFFF0;
    // rom_array[41703] = 32'hFFFFFFF0;
    // rom_array[41704] = 32'hFFFFFFF0;
    // rom_array[41705] = 32'hFFFFFFF1;
    // rom_array[41706] = 32'hFFFFFFF1;
    // rom_array[41707] = 32'hFFFFFFF1;
    // rom_array[41708] = 32'hFFFFFFF1;
    // rom_array[41709] = 32'hFFFFFFF0;
    // rom_array[41710] = 32'hFFFFFFF0;
    // rom_array[41711] = 32'hFFFFFFF0;
    // rom_array[41712] = 32'hFFFFFFF0;
    // rom_array[41713] = 32'hFFFFFFF1;
    // rom_array[41714] = 32'hFFFFFFF1;
    // rom_array[41715] = 32'hFFFFFFF1;
    // rom_array[41716] = 32'hFFFFFFF1;
    // rom_array[41717] = 32'hFFFFFFF0;
    // rom_array[41718] = 32'hFFFFFFF0;
    // rom_array[41719] = 32'hFFFFFFF0;
    // rom_array[41720] = 32'hFFFFFFF0;
    // rom_array[41721] = 32'hFFFFFFF1;
    // rom_array[41722] = 32'hFFFFFFF1;
    // rom_array[41723] = 32'hFFFFFFF1;
    // rom_array[41724] = 32'hFFFFFFF1;
    // rom_array[41725] = 32'hFFFFFFF0;
    // rom_array[41726] = 32'hFFFFFFF0;
    // rom_array[41727] = 32'hFFFFFFF0;
    // rom_array[41728] = 32'hFFFFFFF0;
    // rom_array[41729] = 32'hFFFFFFF1;
    // rom_array[41730] = 32'hFFFFFFF1;
    // rom_array[41731] = 32'hFFFFFFF1;
    // rom_array[41732] = 32'hFFFFFFF1;
    // rom_array[41733] = 32'hFFFFFFF0;
    // rom_array[41734] = 32'hFFFFFFF0;
    // rom_array[41735] = 32'hFFFFFFF0;
    // rom_array[41736] = 32'hFFFFFFF0;
    // rom_array[41737] = 32'hFFFFFFF1;
    // rom_array[41738] = 32'hFFFFFFF1;
    // rom_array[41739] = 32'hFFFFFFF1;
    // rom_array[41740] = 32'hFFFFFFF1;
    // rom_array[41741] = 32'hFFFFFFF0;
    // rom_array[41742] = 32'hFFFFFFF0;
    // rom_array[41743] = 32'hFFFFFFF0;
    // rom_array[41744] = 32'hFFFFFFF0;
    // rom_array[41745] = 32'hFFFFFFF1;
    // rom_array[41746] = 32'hFFFFFFF1;
    // rom_array[41747] = 32'hFFFFFFF1;
    // rom_array[41748] = 32'hFFFFFFF1;
    // rom_array[41749] = 32'hFFFFFFF0;
    // rom_array[41750] = 32'hFFFFFFF0;
    // rom_array[41751] = 32'hFFFFFFF0;
    // rom_array[41752] = 32'hFFFFFFF0;
    // rom_array[41753] = 32'hFFFFFFF1;
    // rom_array[41754] = 32'hFFFFFFF1;
    // rom_array[41755] = 32'hFFFFFFF1;
    // rom_array[41756] = 32'hFFFFFFF1;
    // rom_array[41757] = 32'hFFFFFFF0;
    // rom_array[41758] = 32'hFFFFFFF0;
    // rom_array[41759] = 32'hFFFFFFF0;
    // rom_array[41760] = 32'hFFFFFFF0;
    // rom_array[41761] = 32'hFFFFFFF1;
    // rom_array[41762] = 32'hFFFFFFF1;
    // rom_array[41763] = 32'hFFFFFFF1;
    // rom_array[41764] = 32'hFFFFFFF1;
    // rom_array[41765] = 32'hFFFFFFF0;
    // rom_array[41766] = 32'hFFFFFFF0;
    // rom_array[41767] = 32'hFFFFFFF0;
    // rom_array[41768] = 32'hFFFFFFF0;
    // rom_array[41769] = 32'hFFFFFFF1;
    // rom_array[41770] = 32'hFFFFFFF1;
    // rom_array[41771] = 32'hFFFFFFF1;
    // rom_array[41772] = 32'hFFFFFFF1;
    // rom_array[41773] = 32'hFFFFFFF0;
    // rom_array[41774] = 32'hFFFFFFF0;
    // rom_array[41775] = 32'hFFFFFFF0;
    // rom_array[41776] = 32'hFFFFFFF0;
    // rom_array[41777] = 32'hFFFFFFF1;
    // rom_array[41778] = 32'hFFFFFFF1;
    // rom_array[41779] = 32'hFFFFFFF1;
    // rom_array[41780] = 32'hFFFFFFF1;
    // rom_array[41781] = 32'hFFFFFFF0;
    // rom_array[41782] = 32'hFFFFFFF0;
    // rom_array[41783] = 32'hFFFFFFF0;
    // rom_array[41784] = 32'hFFFFFFF0;
    // rom_array[41785] = 32'hFFFFFFF0;
    // rom_array[41786] = 32'hFFFFFFF0;
    // rom_array[41787] = 32'hFFFFFFF0;
    // rom_array[41788] = 32'hFFFFFFF0;
    // rom_array[41789] = 32'hFFFFFFF1;
    // rom_array[41790] = 32'hFFFFFFF1;
    // rom_array[41791] = 32'hFFFFFFF1;
    // rom_array[41792] = 32'hFFFFFFF1;
    // rom_array[41793] = 32'hFFFFFFF0;
    // rom_array[41794] = 32'hFFFFFFF0;
    // rom_array[41795] = 32'hFFFFFFF0;
    // rom_array[41796] = 32'hFFFFFFF0;
    // rom_array[41797] = 32'hFFFFFFF1;
    // rom_array[41798] = 32'hFFFFFFF1;
    // rom_array[41799] = 32'hFFFFFFF1;
    // rom_array[41800] = 32'hFFFFFFF1;
    // rom_array[41801] = 32'hFFFFFFF0;
    // rom_array[41802] = 32'hFFFFFFF0;
    // rom_array[41803] = 32'hFFFFFFF0;
    // rom_array[41804] = 32'hFFFFFFF0;
    // rom_array[41805] = 32'hFFFFFFF1;
    // rom_array[41806] = 32'hFFFFFFF1;
    // rom_array[41807] = 32'hFFFFFFF1;
    // rom_array[41808] = 32'hFFFFFFF1;
    // rom_array[41809] = 32'hFFFFFFF0;
    // rom_array[41810] = 32'hFFFFFFF0;
    // rom_array[41811] = 32'hFFFFFFF0;
    // rom_array[41812] = 32'hFFFFFFF0;
    // rom_array[41813] = 32'hFFFFFFF1;
    // rom_array[41814] = 32'hFFFFFFF1;
    // rom_array[41815] = 32'hFFFFFFF1;
    // rom_array[41816] = 32'hFFFFFFF1;
    // rom_array[41817] = 32'hFFFFFFF1;
    // rom_array[41818] = 32'hFFFFFFF1;
    // rom_array[41819] = 32'hFFFFFFF1;
    // rom_array[41820] = 32'hFFFFFFF1;
    // rom_array[41821] = 32'hFFFFFFF1;
    // rom_array[41822] = 32'hFFFFFFF1;
    // rom_array[41823] = 32'hFFFFFFF1;
    // rom_array[41824] = 32'hFFFFFFF1;
    // rom_array[41825] = 32'hFFFFFFF1;
    // rom_array[41826] = 32'hFFFFFFF1;
    // rom_array[41827] = 32'hFFFFFFF1;
    // rom_array[41828] = 32'hFFFFFFF1;
    // rom_array[41829] = 32'hFFFFFFF1;
    // rom_array[41830] = 32'hFFFFFFF1;
    // rom_array[41831] = 32'hFFFFFFF1;
    // rom_array[41832] = 32'hFFFFFFF1;
    // rom_array[41833] = 32'hFFFFFFF1;
    // rom_array[41834] = 32'hFFFFFFF1;
    // rom_array[41835] = 32'hFFFFFFF1;
    // rom_array[41836] = 32'hFFFFFFF1;
    // rom_array[41837] = 32'hFFFFFFF1;
    // rom_array[41838] = 32'hFFFFFFF1;
    // rom_array[41839] = 32'hFFFFFFF1;
    // rom_array[41840] = 32'hFFFFFFF1;
    // rom_array[41841] = 32'hFFFFFFF1;
    // rom_array[41842] = 32'hFFFFFFF1;
    // rom_array[41843] = 32'hFFFFFFF1;
    // rom_array[41844] = 32'hFFFFFFF1;
    // rom_array[41845] = 32'hFFFFFFF1;
    // rom_array[41846] = 32'hFFFFFFF1;
    // rom_array[41847] = 32'hFFFFFFF1;
    // rom_array[41848] = 32'hFFFFFFF1;
    // rom_array[41849] = 32'hFFFFFFF1;
    // rom_array[41850] = 32'hFFFFFFF1;
    // rom_array[41851] = 32'hFFFFFFF1;
    // rom_array[41852] = 32'hFFFFFFF1;
    // rom_array[41853] = 32'hFFFFFFF1;
    // rom_array[41854] = 32'hFFFFFFF1;
    // rom_array[41855] = 32'hFFFFFFF1;
    // rom_array[41856] = 32'hFFFFFFF1;
    // rom_array[41857] = 32'hFFFFFFF1;
    // rom_array[41858] = 32'hFFFFFFF1;
    // rom_array[41859] = 32'hFFFFFFF1;
    // rom_array[41860] = 32'hFFFFFFF1;
    // rom_array[41861] = 32'hFFFFFFF1;
    // rom_array[41862] = 32'hFFFFFFF1;
    // rom_array[41863] = 32'hFFFFFFF1;
    // rom_array[41864] = 32'hFFFFFFF1;
    // rom_array[41865] = 32'hFFFFFFF1;
    // rom_array[41866] = 32'hFFFFFFF1;
    // rom_array[41867] = 32'hFFFFFFF1;
    // rom_array[41868] = 32'hFFFFFFF1;
    // rom_array[41869] = 32'hFFFFFFF1;
    // rom_array[41870] = 32'hFFFFFFF1;
    // rom_array[41871] = 32'hFFFFFFF1;
    // rom_array[41872] = 32'hFFFFFFF1;
    // rom_array[41873] = 32'hFFFFFFF1;
    // rom_array[41874] = 32'hFFFFFFF1;
    // rom_array[41875] = 32'hFFFFFFF1;
    // rom_array[41876] = 32'hFFFFFFF1;
    // rom_array[41877] = 32'hFFFFFFF1;
    // rom_array[41878] = 32'hFFFFFFF1;
    // rom_array[41879] = 32'hFFFFFFF1;
    // rom_array[41880] = 32'hFFFFFFF1;
    // rom_array[41881] = 32'hFFFFFFF1;
    // rom_array[41882] = 32'hFFFFFFF1;
    // rom_array[41883] = 32'hFFFFFFF1;
    // rom_array[41884] = 32'hFFFFFFF1;
    // rom_array[41885] = 32'hFFFFFFF0;
    // rom_array[41886] = 32'hFFFFFFF0;
    // rom_array[41887] = 32'hFFFFFFF0;
    // rom_array[41888] = 32'hFFFFFFF0;
    // rom_array[41889] = 32'hFFFFFFF1;
    // rom_array[41890] = 32'hFFFFFFF1;
    // rom_array[41891] = 32'hFFFFFFF1;
    // rom_array[41892] = 32'hFFFFFFF1;
    // rom_array[41893] = 32'hFFFFFFF0;
    // rom_array[41894] = 32'hFFFFFFF0;
    // rom_array[41895] = 32'hFFFFFFF0;
    // rom_array[41896] = 32'hFFFFFFF0;
    // rom_array[41897] = 32'hFFFFFFF1;
    // rom_array[41898] = 32'hFFFFFFF1;
    // rom_array[41899] = 32'hFFFFFFF1;
    // rom_array[41900] = 32'hFFFFFFF1;
    // rom_array[41901] = 32'hFFFFFFF0;
    // rom_array[41902] = 32'hFFFFFFF0;
    // rom_array[41903] = 32'hFFFFFFF0;
    // rom_array[41904] = 32'hFFFFFFF0;
    // rom_array[41905] = 32'hFFFFFFF1;
    // rom_array[41906] = 32'hFFFFFFF1;
    // rom_array[41907] = 32'hFFFFFFF1;
    // rom_array[41908] = 32'hFFFFFFF1;
    // rom_array[41909] = 32'hFFFFFFF0;
    // rom_array[41910] = 32'hFFFFFFF0;
    // rom_array[41911] = 32'hFFFFFFF0;
    // rom_array[41912] = 32'hFFFFFFF0;
    // rom_array[41913] = 32'hFFFFFFF1;
    // rom_array[41914] = 32'hFFFFFFF1;
    // rom_array[41915] = 32'hFFFFFFF1;
    // rom_array[41916] = 32'hFFFFFFF1;
    // rom_array[41917] = 32'hFFFFFFF1;
    // rom_array[41918] = 32'hFFFFFFF1;
    // rom_array[41919] = 32'hFFFFFFF1;
    // rom_array[41920] = 32'hFFFFFFF1;
    // rom_array[41921] = 32'hFFFFFFF1;
    // rom_array[41922] = 32'hFFFFFFF1;
    // rom_array[41923] = 32'hFFFFFFF1;
    // rom_array[41924] = 32'hFFFFFFF1;
    // rom_array[41925] = 32'hFFFFFFF1;
    // rom_array[41926] = 32'hFFFFFFF1;
    // rom_array[41927] = 32'hFFFFFFF1;
    // rom_array[41928] = 32'hFFFFFFF1;
    // rom_array[41929] = 32'hFFFFFFF1;
    // rom_array[41930] = 32'hFFFFFFF1;
    // rom_array[41931] = 32'hFFFFFFF1;
    // rom_array[41932] = 32'hFFFFFFF1;
    // rom_array[41933] = 32'hFFFFFFF1;
    // rom_array[41934] = 32'hFFFFFFF1;
    // rom_array[41935] = 32'hFFFFFFF1;
    // rom_array[41936] = 32'hFFFFFFF1;
    // rom_array[41937] = 32'hFFFFFFF1;
    // rom_array[41938] = 32'hFFFFFFF1;
    // rom_array[41939] = 32'hFFFFFFF1;
    // rom_array[41940] = 32'hFFFFFFF1;
    // rom_array[41941] = 32'hFFFFFFF1;
    // rom_array[41942] = 32'hFFFFFFF1;
    // rom_array[41943] = 32'hFFFFFFF1;
    // rom_array[41944] = 32'hFFFFFFF1;
    // rom_array[41945] = 32'hFFFFFFF1;
    // rom_array[41946] = 32'hFFFFFFF1;
    // rom_array[41947] = 32'hFFFFFFF1;
    // rom_array[41948] = 32'hFFFFFFF1;
    // rom_array[41949] = 32'hFFFFFFF1;
    // rom_array[41950] = 32'hFFFFFFF1;
    // rom_array[41951] = 32'hFFFFFFF1;
    // rom_array[41952] = 32'hFFFFFFF1;
    // rom_array[41953] = 32'hFFFFFFF1;
    // rom_array[41954] = 32'hFFFFFFF1;
    // rom_array[41955] = 32'hFFFFFFF1;
    // rom_array[41956] = 32'hFFFFFFF1;
    // rom_array[41957] = 32'hFFFFFFF1;
    // rom_array[41958] = 32'hFFFFFFF1;
    // rom_array[41959] = 32'hFFFFFFF1;
    // rom_array[41960] = 32'hFFFFFFF1;
    // rom_array[41961] = 32'hFFFFFFF1;
    // rom_array[41962] = 32'hFFFFFFF1;
    // rom_array[41963] = 32'hFFFFFFF1;
    // rom_array[41964] = 32'hFFFFFFF1;
    // rom_array[41965] = 32'hFFFFFFF1;
    // rom_array[41966] = 32'hFFFFFFF1;
    // rom_array[41967] = 32'hFFFFFFF1;
    // rom_array[41968] = 32'hFFFFFFF1;
    // rom_array[41969] = 32'hFFFFFFF1;
    // rom_array[41970] = 32'hFFFFFFF1;
    // rom_array[41971] = 32'hFFFFFFF1;
    // rom_array[41972] = 32'hFFFFFFF1;
    // rom_array[41973] = 32'hFFFFFFF1;
    // rom_array[41974] = 32'hFFFFFFF1;
    // rom_array[41975] = 32'hFFFFFFF1;
    // rom_array[41976] = 32'hFFFFFFF1;
    // rom_array[41977] = 32'hFFFFFFF1;
    // rom_array[41978] = 32'hFFFFFFF1;
    // rom_array[41979] = 32'hFFFFFFF1;
    // rom_array[41980] = 32'hFFFFFFF1;
    // rom_array[41981] = 32'hFFFFFFF0;
    // rom_array[41982] = 32'hFFFFFFF0;
    // rom_array[41983] = 32'hFFFFFFF0;
    // rom_array[41984] = 32'hFFFFFFF0;
    // rom_array[41985] = 32'hFFFFFFF1;
    // rom_array[41986] = 32'hFFFFFFF1;
    // rom_array[41987] = 32'hFFFFFFF1;
    // rom_array[41988] = 32'hFFFFFFF1;
    // rom_array[41989] = 32'hFFFFFFF0;
    // rom_array[41990] = 32'hFFFFFFF0;
    // rom_array[41991] = 32'hFFFFFFF0;
    // rom_array[41992] = 32'hFFFFFFF0;
    // rom_array[41993] = 32'hFFFFFFF1;
    // rom_array[41994] = 32'hFFFFFFF1;
    // rom_array[41995] = 32'hFFFFFFF1;
    // rom_array[41996] = 32'hFFFFFFF1;
    // rom_array[41997] = 32'hFFFFFFF0;
    // rom_array[41998] = 32'hFFFFFFF0;
    // rom_array[41999] = 32'hFFFFFFF0;
    // rom_array[42000] = 32'hFFFFFFF0;
    // rom_array[42001] = 32'hFFFFFFF1;
    // rom_array[42002] = 32'hFFFFFFF1;
    // rom_array[42003] = 32'hFFFFFFF1;
    // rom_array[42004] = 32'hFFFFFFF1;
    // rom_array[42005] = 32'hFFFFFFF0;
    // rom_array[42006] = 32'hFFFFFFF0;
    // rom_array[42007] = 32'hFFFFFFF0;
    // rom_array[42008] = 32'hFFFFFFF0;
    // rom_array[42009] = 32'hFFFFFFF1;
    // rom_array[42010] = 32'hFFFFFFF1;
    // rom_array[42011] = 32'hFFFFFFF1;
    // rom_array[42012] = 32'hFFFFFFF1;
    // rom_array[42013] = 32'hFFFFFFF0;
    // rom_array[42014] = 32'hFFFFFFF0;
    // rom_array[42015] = 32'hFFFFFFF0;
    // rom_array[42016] = 32'hFFFFFFF0;
    // rom_array[42017] = 32'hFFFFFFF1;
    // rom_array[42018] = 32'hFFFFFFF1;
    // rom_array[42019] = 32'hFFFFFFF1;
    // rom_array[42020] = 32'hFFFFFFF1;
    // rom_array[42021] = 32'hFFFFFFF0;
    // rom_array[42022] = 32'hFFFFFFF0;
    // rom_array[42023] = 32'hFFFFFFF0;
    // rom_array[42024] = 32'hFFFFFFF0;
    // rom_array[42025] = 32'hFFFFFFF1;
    // rom_array[42026] = 32'hFFFFFFF1;
    // rom_array[42027] = 32'hFFFFFFF1;
    // rom_array[42028] = 32'hFFFFFFF1;
    // rom_array[42029] = 32'hFFFFFFF0;
    // rom_array[42030] = 32'hFFFFFFF0;
    // rom_array[42031] = 32'hFFFFFFF0;
    // rom_array[42032] = 32'hFFFFFFF0;
    // rom_array[42033] = 32'hFFFFFFF1;
    // rom_array[42034] = 32'hFFFFFFF1;
    // rom_array[42035] = 32'hFFFFFFF1;
    // rom_array[42036] = 32'hFFFFFFF1;
    // rom_array[42037] = 32'hFFFFFFF0;
    // rom_array[42038] = 32'hFFFFFFF0;
    // rom_array[42039] = 32'hFFFFFFF0;
    // rom_array[42040] = 32'hFFFFFFF0;
    // rom_array[42041] = 32'hFFFFFFF1;
    // rom_array[42042] = 32'hFFFFFFF1;
    // rom_array[42043] = 32'hFFFFFFF1;
    // rom_array[42044] = 32'hFFFFFFF1;
    // rom_array[42045] = 32'hFFFFFFF0;
    // rom_array[42046] = 32'hFFFFFFF0;
    // rom_array[42047] = 32'hFFFFFFF0;
    // rom_array[42048] = 32'hFFFFFFF0;
    // rom_array[42049] = 32'hFFFFFFF1;
    // rom_array[42050] = 32'hFFFFFFF1;
    // rom_array[42051] = 32'hFFFFFFF1;
    // rom_array[42052] = 32'hFFFFFFF1;
    // rom_array[42053] = 32'hFFFFFFF0;
    // rom_array[42054] = 32'hFFFFFFF0;
    // rom_array[42055] = 32'hFFFFFFF0;
    // rom_array[42056] = 32'hFFFFFFF0;
    // rom_array[42057] = 32'hFFFFFFF1;
    // rom_array[42058] = 32'hFFFFFFF1;
    // rom_array[42059] = 32'hFFFFFFF1;
    // rom_array[42060] = 32'hFFFFFFF1;
    // rom_array[42061] = 32'hFFFFFFF0;
    // rom_array[42062] = 32'hFFFFFFF0;
    // rom_array[42063] = 32'hFFFFFFF0;
    // rom_array[42064] = 32'hFFFFFFF0;
    // rom_array[42065] = 32'hFFFFFFF1;
    // rom_array[42066] = 32'hFFFFFFF1;
    // rom_array[42067] = 32'hFFFFFFF1;
    // rom_array[42068] = 32'hFFFFFFF1;
    // rom_array[42069] = 32'hFFFFFFF0;
    // rom_array[42070] = 32'hFFFFFFF0;
    // rom_array[42071] = 32'hFFFFFFF0;
    // rom_array[42072] = 32'hFFFFFFF0;
    // rom_array[42073] = 32'hFFFFFFF1;
    // rom_array[42074] = 32'hFFFFFFF1;
    // rom_array[42075] = 32'hFFFFFFF1;
    // rom_array[42076] = 32'hFFFFFFF1;
    // rom_array[42077] = 32'hFFFFFFF0;
    // rom_array[42078] = 32'hFFFFFFF0;
    // rom_array[42079] = 32'hFFFFFFF0;
    // rom_array[42080] = 32'hFFFFFFF0;
    // rom_array[42081] = 32'hFFFFFFF1;
    // rom_array[42082] = 32'hFFFFFFF1;
    // rom_array[42083] = 32'hFFFFFFF1;
    // rom_array[42084] = 32'hFFFFFFF1;
    // rom_array[42085] = 32'hFFFFFFF0;
    // rom_array[42086] = 32'hFFFFFFF0;
    // rom_array[42087] = 32'hFFFFFFF0;
    // rom_array[42088] = 32'hFFFFFFF0;
    // rom_array[42089] = 32'hFFFFFFF1;
    // rom_array[42090] = 32'hFFFFFFF1;
    // rom_array[42091] = 32'hFFFFFFF1;
    // rom_array[42092] = 32'hFFFFFFF1;
    // rom_array[42093] = 32'hFFFFFFF0;
    // rom_array[42094] = 32'hFFFFFFF0;
    // rom_array[42095] = 32'hFFFFFFF0;
    // rom_array[42096] = 32'hFFFFFFF0;
    // rom_array[42097] = 32'hFFFFFFF1;
    // rom_array[42098] = 32'hFFFFFFF1;
    // rom_array[42099] = 32'hFFFFFFF1;
    // rom_array[42100] = 32'hFFFFFFF1;
    // rom_array[42101] = 32'hFFFFFFF0;
    // rom_array[42102] = 32'hFFFFFFF0;
    // rom_array[42103] = 32'hFFFFFFF0;
    // rom_array[42104] = 32'hFFFFFFF0;
    // rom_array[42105] = 32'hFFFFFFF1;
    // rom_array[42106] = 32'hFFFFFFF1;
    // rom_array[42107] = 32'hFFFFFFF1;
    // rom_array[42108] = 32'hFFFFFFF1;
    // rom_array[42109] = 32'hFFFFFFF1;
    // rom_array[42110] = 32'hFFFFFFF1;
    // rom_array[42111] = 32'hFFFFFFF1;
    // rom_array[42112] = 32'hFFFFFFF1;
    // rom_array[42113] = 32'hFFFFFFF1;
    // rom_array[42114] = 32'hFFFFFFF1;
    // rom_array[42115] = 32'hFFFFFFF1;
    // rom_array[42116] = 32'hFFFFFFF1;
    // rom_array[42117] = 32'hFFFFFFF1;
    // rom_array[42118] = 32'hFFFFFFF1;
    // rom_array[42119] = 32'hFFFFFFF1;
    // rom_array[42120] = 32'hFFFFFFF1;
    // rom_array[42121] = 32'hFFFFFFF1;
    // rom_array[42122] = 32'hFFFFFFF1;
    // rom_array[42123] = 32'hFFFFFFF1;
    // rom_array[42124] = 32'hFFFFFFF1;
    // rom_array[42125] = 32'hFFFFFFF1;
    // rom_array[42126] = 32'hFFFFFFF1;
    // rom_array[42127] = 32'hFFFFFFF1;
    // rom_array[42128] = 32'hFFFFFFF1;
    // rom_array[42129] = 32'hFFFFFFF1;
    // rom_array[42130] = 32'hFFFFFFF1;
    // rom_array[42131] = 32'hFFFFFFF1;
    // rom_array[42132] = 32'hFFFFFFF1;
    // rom_array[42133] = 32'hFFFFFFF1;
    // rom_array[42134] = 32'hFFFFFFF1;
    // rom_array[42135] = 32'hFFFFFFF1;
    // rom_array[42136] = 32'hFFFFFFF1;
    // rom_array[42137] = 32'hFFFFFFF1;
    // rom_array[42138] = 32'hFFFFFFF1;
    // rom_array[42139] = 32'hFFFFFFF1;
    // rom_array[42140] = 32'hFFFFFFF1;
    // rom_array[42141] = 32'hFFFFFFF1;
    // rom_array[42142] = 32'hFFFFFFF1;
    // rom_array[42143] = 32'hFFFFFFF1;
    // rom_array[42144] = 32'hFFFFFFF1;
    // rom_array[42145] = 32'hFFFFFFF1;
    // rom_array[42146] = 32'hFFFFFFF1;
    // rom_array[42147] = 32'hFFFFFFF1;
    // rom_array[42148] = 32'hFFFFFFF1;
    // rom_array[42149] = 32'hFFFFFFF1;
    // rom_array[42150] = 32'hFFFFFFF1;
    // rom_array[42151] = 32'hFFFFFFF1;
    // rom_array[42152] = 32'hFFFFFFF1;
    // rom_array[42153] = 32'hFFFFFFF1;
    // rom_array[42154] = 32'hFFFFFFF1;
    // rom_array[42155] = 32'hFFFFFFF1;
    // rom_array[42156] = 32'hFFFFFFF1;
    // rom_array[42157] = 32'hFFFFFFF1;
    // rom_array[42158] = 32'hFFFFFFF1;
    // rom_array[42159] = 32'hFFFFFFF1;
    // rom_array[42160] = 32'hFFFFFFF1;
    // rom_array[42161] = 32'hFFFFFFF1;
    // rom_array[42162] = 32'hFFFFFFF1;
    // rom_array[42163] = 32'hFFFFFFF1;
    // rom_array[42164] = 32'hFFFFFFF1;
    // rom_array[42165] = 32'hFFFFFFF1;
    // rom_array[42166] = 32'hFFFFFFF1;
    // rom_array[42167] = 32'hFFFFFFF1;
    // rom_array[42168] = 32'hFFFFFFF1;
    // rom_array[42169] = 32'hFFFFFFF1;
    // rom_array[42170] = 32'hFFFFFFF1;
    // rom_array[42171] = 32'hFFFFFFF1;
    // rom_array[42172] = 32'hFFFFFFF1;
    // rom_array[42173] = 32'hFFFFFFF0;
    // rom_array[42174] = 32'hFFFFFFF0;
    // rom_array[42175] = 32'hFFFFFFF0;
    // rom_array[42176] = 32'hFFFFFFF0;
    // rom_array[42177] = 32'hFFFFFFF1;
    // rom_array[42178] = 32'hFFFFFFF1;
    // rom_array[42179] = 32'hFFFFFFF1;
    // rom_array[42180] = 32'hFFFFFFF1;
    // rom_array[42181] = 32'hFFFFFFF0;
    // rom_array[42182] = 32'hFFFFFFF0;
    // rom_array[42183] = 32'hFFFFFFF0;
    // rom_array[42184] = 32'hFFFFFFF0;
    // rom_array[42185] = 32'hFFFFFFF1;
    // rom_array[42186] = 32'hFFFFFFF1;
    // rom_array[42187] = 32'hFFFFFFF1;
    // rom_array[42188] = 32'hFFFFFFF1;
    // rom_array[42189] = 32'hFFFFFFF0;
    // rom_array[42190] = 32'hFFFFFFF0;
    // rom_array[42191] = 32'hFFFFFFF0;
    // rom_array[42192] = 32'hFFFFFFF0;
    // rom_array[42193] = 32'hFFFFFFF1;
    // rom_array[42194] = 32'hFFFFFFF1;
    // rom_array[42195] = 32'hFFFFFFF1;
    // rom_array[42196] = 32'hFFFFFFF1;
    // rom_array[42197] = 32'hFFFFFFF0;
    // rom_array[42198] = 32'hFFFFFFF0;
    // rom_array[42199] = 32'hFFFFFFF0;
    // rom_array[42200] = 32'hFFFFFFF0;
    // rom_array[42201] = 32'hFFFFFFF1;
    // rom_array[42202] = 32'hFFFFFFF1;
    // rom_array[42203] = 32'hFFFFFFF1;
    // rom_array[42204] = 32'hFFFFFFF1;
    // rom_array[42205] = 32'hFFFFFFF0;
    // rom_array[42206] = 32'hFFFFFFF0;
    // rom_array[42207] = 32'hFFFFFFF0;
    // rom_array[42208] = 32'hFFFFFFF0;
    // rom_array[42209] = 32'hFFFFFFF1;
    // rom_array[42210] = 32'hFFFFFFF1;
    // rom_array[42211] = 32'hFFFFFFF1;
    // rom_array[42212] = 32'hFFFFFFF1;
    // rom_array[42213] = 32'hFFFFFFF0;
    // rom_array[42214] = 32'hFFFFFFF0;
    // rom_array[42215] = 32'hFFFFFFF0;
    // rom_array[42216] = 32'hFFFFFFF0;
    // rom_array[42217] = 32'hFFFFFFF0;
    // rom_array[42218] = 32'hFFFFFFF0;
    // rom_array[42219] = 32'hFFFFFFF0;
    // rom_array[42220] = 32'hFFFFFFF0;
    // rom_array[42221] = 32'hFFFFFFF1;
    // rom_array[42222] = 32'hFFFFFFF1;
    // rom_array[42223] = 32'hFFFFFFF1;
    // rom_array[42224] = 32'hFFFFFFF1;
    // rom_array[42225] = 32'hFFFFFFF0;
    // rom_array[42226] = 32'hFFFFFFF0;
    // rom_array[42227] = 32'hFFFFFFF0;
    // rom_array[42228] = 32'hFFFFFFF0;
    // rom_array[42229] = 32'hFFFFFFF1;
    // rom_array[42230] = 32'hFFFFFFF1;
    // rom_array[42231] = 32'hFFFFFFF1;
    // rom_array[42232] = 32'hFFFFFFF1;
    // rom_array[42233] = 32'hFFFFFFF0;
    // rom_array[42234] = 32'hFFFFFFF0;
    // rom_array[42235] = 32'hFFFFFFF0;
    // rom_array[42236] = 32'hFFFFFFF0;
    // rom_array[42237] = 32'hFFFFFFF1;
    // rom_array[42238] = 32'hFFFFFFF1;
    // rom_array[42239] = 32'hFFFFFFF1;
    // rom_array[42240] = 32'hFFFFFFF1;
    // rom_array[42241] = 32'hFFFFFFF0;
    // rom_array[42242] = 32'hFFFFFFF0;
    // rom_array[42243] = 32'hFFFFFFF0;
    // rom_array[42244] = 32'hFFFFFFF0;
    // rom_array[42245] = 32'hFFFFFFF1;
    // rom_array[42246] = 32'hFFFFFFF1;
    // rom_array[42247] = 32'hFFFFFFF1;
    // rom_array[42248] = 32'hFFFFFFF1;
    // rom_array[42249] = 32'hFFFFFFF0;
    // rom_array[42250] = 32'hFFFFFFF0;
    // rom_array[42251] = 32'hFFFFFFF0;
    // rom_array[42252] = 32'hFFFFFFF0;
    // rom_array[42253] = 32'hFFFFFFF1;
    // rom_array[42254] = 32'hFFFFFFF1;
    // rom_array[42255] = 32'hFFFFFFF1;
    // rom_array[42256] = 32'hFFFFFFF1;
    // rom_array[42257] = 32'hFFFFFFF0;
    // rom_array[42258] = 32'hFFFFFFF0;
    // rom_array[42259] = 32'hFFFFFFF0;
    // rom_array[42260] = 32'hFFFFFFF0;
    // rom_array[42261] = 32'hFFFFFFF1;
    // rom_array[42262] = 32'hFFFFFFF1;
    // rom_array[42263] = 32'hFFFFFFF1;
    // rom_array[42264] = 32'hFFFFFFF1;
    // rom_array[42265] = 32'hFFFFFFF0;
    // rom_array[42266] = 32'hFFFFFFF0;
    // rom_array[42267] = 32'hFFFFFFF0;
    // rom_array[42268] = 32'hFFFFFFF0;
    // rom_array[42269] = 32'hFFFFFFF1;
    // rom_array[42270] = 32'hFFFFFFF1;
    // rom_array[42271] = 32'hFFFFFFF1;
    // rom_array[42272] = 32'hFFFFFFF1;
    // rom_array[42273] = 32'hFFFFFFF0;
    // rom_array[42274] = 32'hFFFFFFF0;
    // rom_array[42275] = 32'hFFFFFFF0;
    // rom_array[42276] = 32'hFFFFFFF0;
    // rom_array[42277] = 32'hFFFFFFF1;
    // rom_array[42278] = 32'hFFFFFFF1;
    // rom_array[42279] = 32'hFFFFFFF1;
    // rom_array[42280] = 32'hFFFFFFF1;
    // rom_array[42281] = 32'hFFFFFFF0;
    // rom_array[42282] = 32'hFFFFFFF0;
    // rom_array[42283] = 32'hFFFFFFF0;
    // rom_array[42284] = 32'hFFFFFFF0;
    // rom_array[42285] = 32'hFFFFFFF1;
    // rom_array[42286] = 32'hFFFFFFF1;
    // rom_array[42287] = 32'hFFFFFFF1;
    // rom_array[42288] = 32'hFFFFFFF1;
    // rom_array[42289] = 32'hFFFFFFF0;
    // rom_array[42290] = 32'hFFFFFFF0;
    // rom_array[42291] = 32'hFFFFFFF0;
    // rom_array[42292] = 32'hFFFFFFF0;
    // rom_array[42293] = 32'hFFFFFFF1;
    // rom_array[42294] = 32'hFFFFFFF1;
    // rom_array[42295] = 32'hFFFFFFF1;
    // rom_array[42296] = 32'hFFFFFFF1;
    // rom_array[42297] = 32'hFFFFFFF0;
    // rom_array[42298] = 32'hFFFFFFF0;
    // rom_array[42299] = 32'hFFFFFFF0;
    // rom_array[42300] = 32'hFFFFFFF0;
    // rom_array[42301] = 32'hFFFFFFF1;
    // rom_array[42302] = 32'hFFFFFFF1;
    // rom_array[42303] = 32'hFFFFFFF1;
    // rom_array[42304] = 32'hFFFFFFF1;
    // rom_array[42305] = 32'hFFFFFFF0;
    // rom_array[42306] = 32'hFFFFFFF0;
    // rom_array[42307] = 32'hFFFFFFF0;
    // rom_array[42308] = 32'hFFFFFFF0;
    // rom_array[42309] = 32'hFFFFFFF1;
    // rom_array[42310] = 32'hFFFFFFF1;
    // rom_array[42311] = 32'hFFFFFFF1;
    // rom_array[42312] = 32'hFFFFFFF1;
    // rom_array[42313] = 32'hFFFFFFF0;
    // rom_array[42314] = 32'hFFFFFFF0;
    // rom_array[42315] = 32'hFFFFFFF0;
    // rom_array[42316] = 32'hFFFFFFF0;
    // rom_array[42317] = 32'hFFFFFFF1;
    // rom_array[42318] = 32'hFFFFFFF1;
    // rom_array[42319] = 32'hFFFFFFF1;
    // rom_array[42320] = 32'hFFFFFFF1;
    // rom_array[42321] = 32'hFFFFFFF0;
    // rom_array[42322] = 32'hFFFFFFF0;
    // rom_array[42323] = 32'hFFFFFFF0;
    // rom_array[42324] = 32'hFFFFFFF0;
    // rom_array[42325] = 32'hFFFFFFF1;
    // rom_array[42326] = 32'hFFFFFFF1;
    // rom_array[42327] = 32'hFFFFFFF1;
    // rom_array[42328] = 32'hFFFFFFF1;
    // rom_array[42329] = 32'hFFFFFFF0;
    // rom_array[42330] = 32'hFFFFFFF0;
    // rom_array[42331] = 32'hFFFFFFF0;
    // rom_array[42332] = 32'hFFFFFFF0;
    // rom_array[42333] = 32'hFFFFFFF1;
    // rom_array[42334] = 32'hFFFFFFF1;
    // rom_array[42335] = 32'hFFFFFFF1;
    // rom_array[42336] = 32'hFFFFFFF1;
    // rom_array[42337] = 32'hFFFFFFF0;
    // rom_array[42338] = 32'hFFFFFFF0;
    // rom_array[42339] = 32'hFFFFFFF0;
    // rom_array[42340] = 32'hFFFFFFF0;
    // rom_array[42341] = 32'hFFFFFFF1;
    // rom_array[42342] = 32'hFFFFFFF1;
    // rom_array[42343] = 32'hFFFFFFF1;
    // rom_array[42344] = 32'hFFFFFFF1;
    // rom_array[42345] = 32'hFFFFFFF0;
    // rom_array[42346] = 32'hFFFFFFF0;
    // rom_array[42347] = 32'hFFFFFFF0;
    // rom_array[42348] = 32'hFFFFFFF0;
    // rom_array[42349] = 32'hFFFFFFF1;
    // rom_array[42350] = 32'hFFFFFFF1;
    // rom_array[42351] = 32'hFFFFFFF1;
    // rom_array[42352] = 32'hFFFFFFF1;
    // rom_array[42353] = 32'hFFFFFFF0;
    // rom_array[42354] = 32'hFFFFFFF0;
    // rom_array[42355] = 32'hFFFFFFF0;
    // rom_array[42356] = 32'hFFFFFFF0;
    // rom_array[42357] = 32'hFFFFFFF1;
    // rom_array[42358] = 32'hFFFFFFF1;
    // rom_array[42359] = 32'hFFFFFFF1;
    // rom_array[42360] = 32'hFFFFFFF1;
    // rom_array[42361] = 32'hFFFFFFF0;
    // rom_array[42362] = 32'hFFFFFFF0;
    // rom_array[42363] = 32'hFFFFFFF0;
    // rom_array[42364] = 32'hFFFFFFF0;
    // rom_array[42365] = 32'hFFFFFFF1;
    // rom_array[42366] = 32'hFFFFFFF1;
    // rom_array[42367] = 32'hFFFFFFF1;
    // rom_array[42368] = 32'hFFFFFFF1;
    // rom_array[42369] = 32'hFFFFFFF0;
    // rom_array[42370] = 32'hFFFFFFF0;
    // rom_array[42371] = 32'hFFFFFFF0;
    // rom_array[42372] = 32'hFFFFFFF0;
    // rom_array[42373] = 32'hFFFFFFF1;
    // rom_array[42374] = 32'hFFFFFFF1;
    // rom_array[42375] = 32'hFFFFFFF1;
    // rom_array[42376] = 32'hFFFFFFF1;
    // rom_array[42377] = 32'hFFFFFFF0;
    // rom_array[42378] = 32'hFFFFFFF0;
    // rom_array[42379] = 32'hFFFFFFF0;
    // rom_array[42380] = 32'hFFFFFFF0;
    // rom_array[42381] = 32'hFFFFFFF1;
    // rom_array[42382] = 32'hFFFFFFF1;
    // rom_array[42383] = 32'hFFFFFFF1;
    // rom_array[42384] = 32'hFFFFFFF1;
    // rom_array[42385] = 32'hFFFFFFF0;
    // rom_array[42386] = 32'hFFFFFFF0;
    // rom_array[42387] = 32'hFFFFFFF0;
    // rom_array[42388] = 32'hFFFFFFF0;
    // rom_array[42389] = 32'hFFFFFFF1;
    // rom_array[42390] = 32'hFFFFFFF1;
    // rom_array[42391] = 32'hFFFFFFF1;
    // rom_array[42392] = 32'hFFFFFFF1;
    // rom_array[42393] = 32'hFFFFFFF1;
    // rom_array[42394] = 32'hFFFFFFF1;
    // rom_array[42395] = 32'hFFFFFFF1;
    // rom_array[42396] = 32'hFFFFFFF1;
    // rom_array[42397] = 32'hFFFFFFF1;
    // rom_array[42398] = 32'hFFFFFFF1;
    // rom_array[42399] = 32'hFFFFFFF1;
    // rom_array[42400] = 32'hFFFFFFF1;
    // rom_array[42401] = 32'hFFFFFFF1;
    // rom_array[42402] = 32'hFFFFFFF1;
    // rom_array[42403] = 32'hFFFFFFF1;
    // rom_array[42404] = 32'hFFFFFFF1;
    // rom_array[42405] = 32'hFFFFFFF1;
    // rom_array[42406] = 32'hFFFFFFF1;
    // rom_array[42407] = 32'hFFFFFFF1;
    // rom_array[42408] = 32'hFFFFFFF1;
    // rom_array[42409] = 32'hFFFFFFF1;
    // rom_array[42410] = 32'hFFFFFFF1;
    // rom_array[42411] = 32'hFFFFFFF1;
    // rom_array[42412] = 32'hFFFFFFF1;
    // rom_array[42413] = 32'hFFFFFFF1;
    // rom_array[42414] = 32'hFFFFFFF1;
    // rom_array[42415] = 32'hFFFFFFF1;
    // rom_array[42416] = 32'hFFFFFFF1;
    // rom_array[42417] = 32'hFFFFFFF1;
    // rom_array[42418] = 32'hFFFFFFF1;
    // rom_array[42419] = 32'hFFFFFFF1;
    // rom_array[42420] = 32'hFFFFFFF1;
    // rom_array[42421] = 32'hFFFFFFF1;
    // rom_array[42422] = 32'hFFFFFFF1;
    // rom_array[42423] = 32'hFFFFFFF1;
    // rom_array[42424] = 32'hFFFFFFF1;
    // rom_array[42425] = 32'hFFFFFFF1;
    // rom_array[42426] = 32'hFFFFFFF1;
    // rom_array[42427] = 32'hFFFFFFF1;
    // rom_array[42428] = 32'hFFFFFFF1;
    // rom_array[42429] = 32'hFFFFFFF1;
    // rom_array[42430] = 32'hFFFFFFF1;
    // rom_array[42431] = 32'hFFFFFFF1;
    // rom_array[42432] = 32'hFFFFFFF1;
    // rom_array[42433] = 32'hFFFFFFF1;
    // rom_array[42434] = 32'hFFFFFFF1;
    // rom_array[42435] = 32'hFFFFFFF1;
    // rom_array[42436] = 32'hFFFFFFF1;
    // rom_array[42437] = 32'hFFFFFFF1;
    // rom_array[42438] = 32'hFFFFFFF1;
    // rom_array[42439] = 32'hFFFFFFF1;
    // rom_array[42440] = 32'hFFFFFFF1;
    // rom_array[42441] = 32'hFFFFFFF1;
    // rom_array[42442] = 32'hFFFFFFF1;
    // rom_array[42443] = 32'hFFFFFFF1;
    // rom_array[42444] = 32'hFFFFFFF1;
    // rom_array[42445] = 32'hFFFFFFF0;
    // rom_array[42446] = 32'hFFFFFFF0;
    // rom_array[42447] = 32'hFFFFFFF0;
    // rom_array[42448] = 32'hFFFFFFF0;
    // rom_array[42449] = 32'hFFFFFFF1;
    // rom_array[42450] = 32'hFFFFFFF1;
    // rom_array[42451] = 32'hFFFFFFF1;
    // rom_array[42452] = 32'hFFFFFFF1;
    // rom_array[42453] = 32'hFFFFFFF0;
    // rom_array[42454] = 32'hFFFFFFF0;
    // rom_array[42455] = 32'hFFFFFFF0;
    // rom_array[42456] = 32'hFFFFFFF0;
    // rom_array[42457] = 32'hFFFFFFF1;
    // rom_array[42458] = 32'hFFFFFFF1;
    // rom_array[42459] = 32'hFFFFFFF1;
    // rom_array[42460] = 32'hFFFFFFF1;
    // rom_array[42461] = 32'hFFFFFFF0;
    // rom_array[42462] = 32'hFFFFFFF0;
    // rom_array[42463] = 32'hFFFFFFF0;
    // rom_array[42464] = 32'hFFFFFFF0;
    // rom_array[42465] = 32'hFFFFFFF1;
    // rom_array[42466] = 32'hFFFFFFF1;
    // rom_array[42467] = 32'hFFFFFFF1;
    // rom_array[42468] = 32'hFFFFFFF1;
    // rom_array[42469] = 32'hFFFFFFF0;
    // rom_array[42470] = 32'hFFFFFFF0;
    // rom_array[42471] = 32'hFFFFFFF0;
    // rom_array[42472] = 32'hFFFFFFF0;
    // rom_array[42473] = 32'hFFFFFFF1;
    // rom_array[42474] = 32'hFFFFFFF1;
    // rom_array[42475] = 32'hFFFFFFF1;
    // rom_array[42476] = 32'hFFFFFFF1;
    // rom_array[42477] = 32'hFFFFFFF0;
    // rom_array[42478] = 32'hFFFFFFF0;
    // rom_array[42479] = 32'hFFFFFFF0;
    // rom_array[42480] = 32'hFFFFFFF0;
    // rom_array[42481] = 32'hFFFFFFF1;
    // rom_array[42482] = 32'hFFFFFFF1;
    // rom_array[42483] = 32'hFFFFFFF1;
    // rom_array[42484] = 32'hFFFFFFF1;
    // rom_array[42485] = 32'hFFFFFFF0;
    // rom_array[42486] = 32'hFFFFFFF0;
    // rom_array[42487] = 32'hFFFFFFF0;
    // rom_array[42488] = 32'hFFFFFFF0;
    // rom_array[42489] = 32'hFFFFFFF1;
    // rom_array[42490] = 32'hFFFFFFF1;
    // rom_array[42491] = 32'hFFFFFFF1;
    // rom_array[42492] = 32'hFFFFFFF1;
    // rom_array[42493] = 32'hFFFFFFF0;
    // rom_array[42494] = 32'hFFFFFFF0;
    // rom_array[42495] = 32'hFFFFFFF0;
    // rom_array[42496] = 32'hFFFFFFF0;
    // rom_array[42497] = 32'hFFFFFFF1;
    // rom_array[42498] = 32'hFFFFFFF1;
    // rom_array[42499] = 32'hFFFFFFF1;
    // rom_array[42500] = 32'hFFFFFFF1;
    // rom_array[42501] = 32'hFFFFFFF0;
    // rom_array[42502] = 32'hFFFFFFF0;
    // rom_array[42503] = 32'hFFFFFFF0;
    // rom_array[42504] = 32'hFFFFFFF0;
    // rom_array[42505] = 32'hFFFFFFF1;
    // rom_array[42506] = 32'hFFFFFFF1;
    // rom_array[42507] = 32'hFFFFFFF1;
    // rom_array[42508] = 32'hFFFFFFF1;
    // rom_array[42509] = 32'hFFFFFFF0;
    // rom_array[42510] = 32'hFFFFFFF0;
    // rom_array[42511] = 32'hFFFFFFF0;
    // rom_array[42512] = 32'hFFFFFFF0;
    // rom_array[42513] = 32'hFFFFFFF1;
    // rom_array[42514] = 32'hFFFFFFF1;
    // rom_array[42515] = 32'hFFFFFFF1;
    // rom_array[42516] = 32'hFFFFFFF1;
    // rom_array[42517] = 32'hFFFFFFF0;
    // rom_array[42518] = 32'hFFFFFFF0;
    // rom_array[42519] = 32'hFFFFFFF0;
    // rom_array[42520] = 32'hFFFFFFF0;
    // rom_array[42521] = 32'hFFFFFFF1;
    // rom_array[42522] = 32'hFFFFFFF1;
    // rom_array[42523] = 32'hFFFFFFF1;
    // rom_array[42524] = 32'hFFFFFFF1;
    // rom_array[42525] = 32'hFFFFFFF0;
    // rom_array[42526] = 32'hFFFFFFF0;
    // rom_array[42527] = 32'hFFFFFFF0;
    // rom_array[42528] = 32'hFFFFFFF0;
    // rom_array[42529] = 32'hFFFFFFF1;
    // rom_array[42530] = 32'hFFFFFFF1;
    // rom_array[42531] = 32'hFFFFFFF1;
    // rom_array[42532] = 32'hFFFFFFF1;
    // rom_array[42533] = 32'hFFFFFFF0;
    // rom_array[42534] = 32'hFFFFFFF0;
    // rom_array[42535] = 32'hFFFFFFF0;
    // rom_array[42536] = 32'hFFFFFFF0;
    // rom_array[42537] = 32'hFFFFFFF1;
    // rom_array[42538] = 32'hFFFFFFF1;
    // rom_array[42539] = 32'hFFFFFFF1;
    // rom_array[42540] = 32'hFFFFFFF1;
    // rom_array[42541] = 32'hFFFFFFF0;
    // rom_array[42542] = 32'hFFFFFFF0;
    // rom_array[42543] = 32'hFFFFFFF0;
    // rom_array[42544] = 32'hFFFFFFF0;
    // rom_array[42545] = 32'hFFFFFFF1;
    // rom_array[42546] = 32'hFFFFFFF1;
    // rom_array[42547] = 32'hFFFFFFF1;
    // rom_array[42548] = 32'hFFFFFFF1;
    // rom_array[42549] = 32'hFFFFFFF0;
    // rom_array[42550] = 32'hFFFFFFF0;
    // rom_array[42551] = 32'hFFFFFFF0;
    // rom_array[42552] = 32'hFFFFFFF0;
    // rom_array[42553] = 32'hFFFFFFF1;
    // rom_array[42554] = 32'hFFFFFFF1;
    // rom_array[42555] = 32'hFFFFFFF1;
    // rom_array[42556] = 32'hFFFFFFF1;
    // rom_array[42557] = 32'hFFFFFFF0;
    // rom_array[42558] = 32'hFFFFFFF0;
    // rom_array[42559] = 32'hFFFFFFF0;
    // rom_array[42560] = 32'hFFFFFFF0;
    // rom_array[42561] = 32'hFFFFFFF1;
    // rom_array[42562] = 32'hFFFFFFF1;
    // rom_array[42563] = 32'hFFFFFFF1;
    // rom_array[42564] = 32'hFFFFFFF1;
    // rom_array[42565] = 32'hFFFFFFF0;
    // rom_array[42566] = 32'hFFFFFFF0;
    // rom_array[42567] = 32'hFFFFFFF0;
    // rom_array[42568] = 32'hFFFFFFF0;
    // rom_array[42569] = 32'hFFFFFFF1;
    // rom_array[42570] = 32'hFFFFFFF1;
    // rom_array[42571] = 32'hFFFFFFF1;
    // rom_array[42572] = 32'hFFFFFFF1;
    // rom_array[42573] = 32'hFFFFFFF0;
    // rom_array[42574] = 32'hFFFFFFF0;
    // rom_array[42575] = 32'hFFFFFFF0;
    // rom_array[42576] = 32'hFFFFFFF0;
    // rom_array[42577] = 32'hFFFFFFF1;
    // rom_array[42578] = 32'hFFFFFFF1;
    // rom_array[42579] = 32'hFFFFFFF1;
    // rom_array[42580] = 32'hFFFFFFF1;
    // rom_array[42581] = 32'hFFFFFFF0;
    // rom_array[42582] = 32'hFFFFFFF0;
    // rom_array[42583] = 32'hFFFFFFF0;
    // rom_array[42584] = 32'hFFFFFFF0;
    // rom_array[42585] = 32'hFFFFFFF1;
    // rom_array[42586] = 32'hFFFFFFF1;
    // rom_array[42587] = 32'hFFFFFFF1;
    // rom_array[42588] = 32'hFFFFFFF1;
    // rom_array[42589] = 32'hFFFFFFF0;
    // rom_array[42590] = 32'hFFFFFFF0;
    // rom_array[42591] = 32'hFFFFFFF0;
    // rom_array[42592] = 32'hFFFFFFF0;
    // rom_array[42593] = 32'hFFFFFFF1;
    // rom_array[42594] = 32'hFFFFFFF1;
    // rom_array[42595] = 32'hFFFFFFF1;
    // rom_array[42596] = 32'hFFFFFFF1;
    // rom_array[42597] = 32'hFFFFFFF0;
    // rom_array[42598] = 32'hFFFFFFF0;
    // rom_array[42599] = 32'hFFFFFFF0;
    // rom_array[42600] = 32'hFFFFFFF0;
    // rom_array[42601] = 32'hFFFFFFF1;
    // rom_array[42602] = 32'hFFFFFFF1;
    // rom_array[42603] = 32'hFFFFFFF1;
    // rom_array[42604] = 32'hFFFFFFF1;
    // rom_array[42605] = 32'hFFFFFFF0;
    // rom_array[42606] = 32'hFFFFFFF0;
    // rom_array[42607] = 32'hFFFFFFF0;
    // rom_array[42608] = 32'hFFFFFFF0;
    // rom_array[42609] = 32'hFFFFFFF1;
    // rom_array[42610] = 32'hFFFFFFF1;
    // rom_array[42611] = 32'hFFFFFFF1;
    // rom_array[42612] = 32'hFFFFFFF1;
    // rom_array[42613] = 32'hFFFFFFF0;
    // rom_array[42614] = 32'hFFFFFFF0;
    // rom_array[42615] = 32'hFFFFFFF0;
    // rom_array[42616] = 32'hFFFFFFF0;
    // rom_array[42617] = 32'hFFFFFFF1;
    // rom_array[42618] = 32'hFFFFFFF1;
    // rom_array[42619] = 32'hFFFFFFF1;
    // rom_array[42620] = 32'hFFFFFFF1;
    // rom_array[42621] = 32'hFFFFFFF0;
    // rom_array[42622] = 32'hFFFFFFF0;
    // rom_array[42623] = 32'hFFFFFFF0;
    // rom_array[42624] = 32'hFFFFFFF0;
    // rom_array[42625] = 32'hFFFFFFF1;
    // rom_array[42626] = 32'hFFFFFFF1;
    // rom_array[42627] = 32'hFFFFFFF1;
    // rom_array[42628] = 32'hFFFFFFF1;
    // rom_array[42629] = 32'hFFFFFFF0;
    // rom_array[42630] = 32'hFFFFFFF0;
    // rom_array[42631] = 32'hFFFFFFF0;
    // rom_array[42632] = 32'hFFFFFFF0;
    // rom_array[42633] = 32'hFFFFFFF1;
    // rom_array[42634] = 32'hFFFFFFF1;
    // rom_array[42635] = 32'hFFFFFFF1;
    // rom_array[42636] = 32'hFFFFFFF1;
    // rom_array[42637] = 32'hFFFFFFF0;
    // rom_array[42638] = 32'hFFFFFFF0;
    // rom_array[42639] = 32'hFFFFFFF0;
    // rom_array[42640] = 32'hFFFFFFF0;
    // rom_array[42641] = 32'hFFFFFFF1;
    // rom_array[42642] = 32'hFFFFFFF1;
    // rom_array[42643] = 32'hFFFFFFF1;
    // rom_array[42644] = 32'hFFFFFFF1;
    // rom_array[42645] = 32'hFFFFFFF0;
    // rom_array[42646] = 32'hFFFFFFF0;
    // rom_array[42647] = 32'hFFFFFFF0;
    // rom_array[42648] = 32'hFFFFFFF0;
    // rom_array[42649] = 32'hFFFFFFF0;
    // rom_array[42650] = 32'hFFFFFFF0;
    // rom_array[42651] = 32'hFFFFFFF1;
    // rom_array[42652] = 32'hFFFFFFF1;
    // rom_array[42653] = 32'hFFFFFFF0;
    // rom_array[42654] = 32'hFFFFFFF0;
    // rom_array[42655] = 32'hFFFFFFF0;
    // rom_array[42656] = 32'hFFFFFFF0;
    // rom_array[42657] = 32'hFFFFFFF0;
    // rom_array[42658] = 32'hFFFFFFF0;
    // rom_array[42659] = 32'hFFFFFFF1;
    // rom_array[42660] = 32'hFFFFFFF1;
    // rom_array[42661] = 32'hFFFFFFF0;
    // rom_array[42662] = 32'hFFFFFFF0;
    // rom_array[42663] = 32'hFFFFFFF0;
    // rom_array[42664] = 32'hFFFFFFF0;
    // rom_array[42665] = 32'hFFFFFFF1;
    // rom_array[42666] = 32'hFFFFFFF1;
    // rom_array[42667] = 32'hFFFFFFF1;
    // rom_array[42668] = 32'hFFFFFFF1;
    // rom_array[42669] = 32'hFFFFFFF0;
    // rom_array[42670] = 32'hFFFFFFF0;
    // rom_array[42671] = 32'hFFFFFFF0;
    // rom_array[42672] = 32'hFFFFFFF0;
    // rom_array[42673] = 32'hFFFFFFF1;
    // rom_array[42674] = 32'hFFFFFFF1;
    // rom_array[42675] = 32'hFFFFFFF1;
    // rom_array[42676] = 32'hFFFFFFF1;
    // rom_array[42677] = 32'hFFFFFFF0;
    // rom_array[42678] = 32'hFFFFFFF0;
    // rom_array[42679] = 32'hFFFFFFF0;
    // rom_array[42680] = 32'hFFFFFFF0;
    // rom_array[42681] = 32'hFFFFFFF1;
    // rom_array[42682] = 32'hFFFFFFF1;
    // rom_array[42683] = 32'hFFFFFFF1;
    // rom_array[42684] = 32'hFFFFFFF1;
    // rom_array[42685] = 32'hFFFFFFF0;
    // rom_array[42686] = 32'hFFFFFFF0;
    // rom_array[42687] = 32'hFFFFFFF0;
    // rom_array[42688] = 32'hFFFFFFF0;
    // rom_array[42689] = 32'hFFFFFFF1;
    // rom_array[42690] = 32'hFFFFFFF1;
    // rom_array[42691] = 32'hFFFFFFF1;
    // rom_array[42692] = 32'hFFFFFFF1;
    // rom_array[42693] = 32'hFFFFFFF0;
    // rom_array[42694] = 32'hFFFFFFF0;
    // rom_array[42695] = 32'hFFFFFFF0;
    // rom_array[42696] = 32'hFFFFFFF0;
    // rom_array[42697] = 32'hFFFFFFF1;
    // rom_array[42698] = 32'hFFFFFFF1;
    // rom_array[42699] = 32'hFFFFFFF1;
    // rom_array[42700] = 32'hFFFFFFF1;
    // rom_array[42701] = 32'hFFFFFFF0;
    // rom_array[42702] = 32'hFFFFFFF0;
    // rom_array[42703] = 32'hFFFFFFF0;
    // rom_array[42704] = 32'hFFFFFFF0;
    // rom_array[42705] = 32'hFFFFFFF1;
    // rom_array[42706] = 32'hFFFFFFF1;
    // rom_array[42707] = 32'hFFFFFFF1;
    // rom_array[42708] = 32'hFFFFFFF1;
    // rom_array[42709] = 32'hFFFFFFF0;
    // rom_array[42710] = 32'hFFFFFFF0;
    // rom_array[42711] = 32'hFFFFFFF0;
    // rom_array[42712] = 32'hFFFFFFF0;
    // rom_array[42713] = 32'hFFFFFFF1;
    // rom_array[42714] = 32'hFFFFFFF1;
    // rom_array[42715] = 32'hFFFFFFF1;
    // rom_array[42716] = 32'hFFFFFFF1;
    // rom_array[42717] = 32'hFFFFFFF0;
    // rom_array[42718] = 32'hFFFFFFF0;
    // rom_array[42719] = 32'hFFFFFFF0;
    // rom_array[42720] = 32'hFFFFFFF0;
    // rom_array[42721] = 32'hFFFFFFF1;
    // rom_array[42722] = 32'hFFFFFFF1;
    // rom_array[42723] = 32'hFFFFFFF1;
    // rom_array[42724] = 32'hFFFFFFF1;
    // rom_array[42725] = 32'hFFFFFFF0;
    // rom_array[42726] = 32'hFFFFFFF0;
    // rom_array[42727] = 32'hFFFFFFF0;
    // rom_array[42728] = 32'hFFFFFFF0;
    // rom_array[42729] = 32'hFFFFFFF0;
    // rom_array[42730] = 32'hFFFFFFF0;
    // rom_array[42731] = 32'hFFFFFFF0;
    // rom_array[42732] = 32'hFFFFFFF0;
    // rom_array[42733] = 32'hFFFFFFF1;
    // rom_array[42734] = 32'hFFFFFFF1;
    // rom_array[42735] = 32'hFFFFFFF1;
    // rom_array[42736] = 32'hFFFFFFF1;
    // rom_array[42737] = 32'hFFFFFFF0;
    // rom_array[42738] = 32'hFFFFFFF0;
    // rom_array[42739] = 32'hFFFFFFF0;
    // rom_array[42740] = 32'hFFFFFFF0;
    // rom_array[42741] = 32'hFFFFFFF1;
    // rom_array[42742] = 32'hFFFFFFF1;
    // rom_array[42743] = 32'hFFFFFFF1;
    // rom_array[42744] = 32'hFFFFFFF1;
    // rom_array[42745] = 32'hFFFFFFF0;
    // rom_array[42746] = 32'hFFFFFFF0;
    // rom_array[42747] = 32'hFFFFFFF0;
    // rom_array[42748] = 32'hFFFFFFF0;
    // rom_array[42749] = 32'hFFFFFFF1;
    // rom_array[42750] = 32'hFFFFFFF1;
    // rom_array[42751] = 32'hFFFFFFF1;
    // rom_array[42752] = 32'hFFFFFFF1;
    // rom_array[42753] = 32'hFFFFFFF0;
    // rom_array[42754] = 32'hFFFFFFF0;
    // rom_array[42755] = 32'hFFFFFFF0;
    // rom_array[42756] = 32'hFFFFFFF0;
    // rom_array[42757] = 32'hFFFFFFF1;
    // rom_array[42758] = 32'hFFFFFFF1;
    // rom_array[42759] = 32'hFFFFFFF1;
    // rom_array[42760] = 32'hFFFFFFF1;
    // rom_array[42761] = 32'hFFFFFFF0;
    // rom_array[42762] = 32'hFFFFFFF0;
    // rom_array[42763] = 32'hFFFFFFF0;
    // rom_array[42764] = 32'hFFFFFFF0;
    // rom_array[42765] = 32'hFFFFFFF1;
    // rom_array[42766] = 32'hFFFFFFF1;
    // rom_array[42767] = 32'hFFFFFFF1;
    // rom_array[42768] = 32'hFFFFFFF1;
    // rom_array[42769] = 32'hFFFFFFF0;
    // rom_array[42770] = 32'hFFFFFFF0;
    // rom_array[42771] = 32'hFFFFFFF0;
    // rom_array[42772] = 32'hFFFFFFF0;
    // rom_array[42773] = 32'hFFFFFFF1;
    // rom_array[42774] = 32'hFFFFFFF1;
    // rom_array[42775] = 32'hFFFFFFF1;
    // rom_array[42776] = 32'hFFFFFFF1;
    // rom_array[42777] = 32'hFFFFFFF0;
    // rom_array[42778] = 32'hFFFFFFF0;
    // rom_array[42779] = 32'hFFFFFFF0;
    // rom_array[42780] = 32'hFFFFFFF0;
    // rom_array[42781] = 32'hFFFFFFF1;
    // rom_array[42782] = 32'hFFFFFFF1;
    // rom_array[42783] = 32'hFFFFFFF1;
    // rom_array[42784] = 32'hFFFFFFF1;
    // rom_array[42785] = 32'hFFFFFFF0;
    // rom_array[42786] = 32'hFFFFFFF0;
    // rom_array[42787] = 32'hFFFFFFF0;
    // rom_array[42788] = 32'hFFFFFFF0;
    // rom_array[42789] = 32'hFFFFFFF1;
    // rom_array[42790] = 32'hFFFFFFF1;
    // rom_array[42791] = 32'hFFFFFFF1;
    // rom_array[42792] = 32'hFFFFFFF1;
    // rom_array[42793] = 32'hFFFFFFF0;
    // rom_array[42794] = 32'hFFFFFFF0;
    // rom_array[42795] = 32'hFFFFFFF0;
    // rom_array[42796] = 32'hFFFFFFF0;
    // rom_array[42797] = 32'hFFFFFFF1;
    // rom_array[42798] = 32'hFFFFFFF1;
    // rom_array[42799] = 32'hFFFFFFF1;
    // rom_array[42800] = 32'hFFFFFFF1;
    // rom_array[42801] = 32'hFFFFFFF0;
    // rom_array[42802] = 32'hFFFFFFF0;
    // rom_array[42803] = 32'hFFFFFFF0;
    // rom_array[42804] = 32'hFFFFFFF0;
    // rom_array[42805] = 32'hFFFFFFF1;
    // rom_array[42806] = 32'hFFFFFFF1;
    // rom_array[42807] = 32'hFFFFFFF1;
    // rom_array[42808] = 32'hFFFFFFF1;
    // rom_array[42809] = 32'hFFFFFFF0;
    // rom_array[42810] = 32'hFFFFFFF0;
    // rom_array[42811] = 32'hFFFFFFF0;
    // rom_array[42812] = 32'hFFFFFFF0;
    // rom_array[42813] = 32'hFFFFFFF1;
    // rom_array[42814] = 32'hFFFFFFF1;
    // rom_array[42815] = 32'hFFFFFFF1;
    // rom_array[42816] = 32'hFFFFFFF1;
    // rom_array[42817] = 32'hFFFFFFF0;
    // rom_array[42818] = 32'hFFFFFFF0;
    // rom_array[42819] = 32'hFFFFFFF0;
    // rom_array[42820] = 32'hFFFFFFF0;
    // rom_array[42821] = 32'hFFFFFFF1;
    // rom_array[42822] = 32'hFFFFFFF1;
    // rom_array[42823] = 32'hFFFFFFF1;
    // rom_array[42824] = 32'hFFFFFFF1;
    // rom_array[42825] = 32'hFFFFFFF0;
    // rom_array[42826] = 32'hFFFFFFF0;
    // rom_array[42827] = 32'hFFFFFFF0;
    // rom_array[42828] = 32'hFFFFFFF0;
    // rom_array[42829] = 32'hFFFFFFF1;
    // rom_array[42830] = 32'hFFFFFFF1;
    // rom_array[42831] = 32'hFFFFFFF1;
    // rom_array[42832] = 32'hFFFFFFF1;
    // rom_array[42833] = 32'hFFFFFFF0;
    // rom_array[42834] = 32'hFFFFFFF0;
    // rom_array[42835] = 32'hFFFFFFF0;
    // rom_array[42836] = 32'hFFFFFFF0;
    // rom_array[42837] = 32'hFFFFFFF1;
    // rom_array[42838] = 32'hFFFFFFF1;
    // rom_array[42839] = 32'hFFFFFFF1;
    // rom_array[42840] = 32'hFFFFFFF1;
    // rom_array[42841] = 32'hFFFFFFF0;
    // rom_array[42842] = 32'hFFFFFFF0;
    // rom_array[42843] = 32'hFFFFFFF0;
    // rom_array[42844] = 32'hFFFFFFF0;
    // rom_array[42845] = 32'hFFFFFFF1;
    // rom_array[42846] = 32'hFFFFFFF1;
    // rom_array[42847] = 32'hFFFFFFF1;
    // rom_array[42848] = 32'hFFFFFFF1;
    // rom_array[42849] = 32'hFFFFFFF0;
    // rom_array[42850] = 32'hFFFFFFF0;
    // rom_array[42851] = 32'hFFFFFFF0;
    // rom_array[42852] = 32'hFFFFFFF0;
    // rom_array[42853] = 32'hFFFFFFF1;
    // rom_array[42854] = 32'hFFFFFFF1;
    // rom_array[42855] = 32'hFFFFFFF1;
    // rom_array[42856] = 32'hFFFFFFF1;
    // rom_array[42857] = 32'hFFFFFFF1;
    // rom_array[42858] = 32'hFFFFFFF1;
    // rom_array[42859] = 32'hFFFFFFF1;
    // rom_array[42860] = 32'hFFFFFFF1;
    // rom_array[42861] = 32'hFFFFFFF1;
    // rom_array[42862] = 32'hFFFFFFF1;
    // rom_array[42863] = 32'hFFFFFFF1;
    // rom_array[42864] = 32'hFFFFFFF1;
    // rom_array[42865] = 32'hFFFFFFF1;
    // rom_array[42866] = 32'hFFFFFFF1;
    // rom_array[42867] = 32'hFFFFFFF1;
    // rom_array[42868] = 32'hFFFFFFF1;
    // rom_array[42869] = 32'hFFFFFFF1;
    // rom_array[42870] = 32'hFFFFFFF1;
    // rom_array[42871] = 32'hFFFFFFF1;
    // rom_array[42872] = 32'hFFFFFFF1;
    // rom_array[42873] = 32'hFFFFFFF1;
    // rom_array[42874] = 32'hFFFFFFF1;
    // rom_array[42875] = 32'hFFFFFFF1;
    // rom_array[42876] = 32'hFFFFFFF1;
    // rom_array[42877] = 32'hFFFFFFF0;
    // rom_array[42878] = 32'hFFFFFFF0;
    // rom_array[42879] = 32'hFFFFFFF0;
    // rom_array[42880] = 32'hFFFFFFF0;
    // rom_array[42881] = 32'hFFFFFFF1;
    // rom_array[42882] = 32'hFFFFFFF1;
    // rom_array[42883] = 32'hFFFFFFF1;
    // rom_array[42884] = 32'hFFFFFFF1;
    // rom_array[42885] = 32'hFFFFFFF0;
    // rom_array[42886] = 32'hFFFFFFF0;
    // rom_array[42887] = 32'hFFFFFFF0;
    // rom_array[42888] = 32'hFFFFFFF0;
    // rom_array[42889] = 32'hFFFFFFF1;
    // rom_array[42890] = 32'hFFFFFFF1;
    // rom_array[42891] = 32'hFFFFFFF1;
    // rom_array[42892] = 32'hFFFFFFF1;
    // rom_array[42893] = 32'hFFFFFFF1;
    // rom_array[42894] = 32'hFFFFFFF1;
    // rom_array[42895] = 32'hFFFFFFF1;
    // rom_array[42896] = 32'hFFFFFFF1;
    // rom_array[42897] = 32'hFFFFFFF1;
    // rom_array[42898] = 32'hFFFFFFF1;
    // rom_array[42899] = 32'hFFFFFFF1;
    // rom_array[42900] = 32'hFFFFFFF1;
    // rom_array[42901] = 32'hFFFFFFF1;
    // rom_array[42902] = 32'hFFFFFFF1;
    // rom_array[42903] = 32'hFFFFFFF1;
    // rom_array[42904] = 32'hFFFFFFF1;
    // rom_array[42905] = 32'hFFFFFFF1;
    // rom_array[42906] = 32'hFFFFFFF1;
    // rom_array[42907] = 32'hFFFFFFF1;
    // rom_array[42908] = 32'hFFFFFFF1;
    // rom_array[42909] = 32'hFFFFFFF0;
    // rom_array[42910] = 32'hFFFFFFF0;
    // rom_array[42911] = 32'hFFFFFFF0;
    // rom_array[42912] = 32'hFFFFFFF0;
    // rom_array[42913] = 32'hFFFFFFF1;
    // rom_array[42914] = 32'hFFFFFFF1;
    // rom_array[42915] = 32'hFFFFFFF1;
    // rom_array[42916] = 32'hFFFFFFF1;
    // rom_array[42917] = 32'hFFFFFFF0;
    // rom_array[42918] = 32'hFFFFFFF0;
    // rom_array[42919] = 32'hFFFFFFF0;
    // rom_array[42920] = 32'hFFFFFFF0;
    // rom_array[42921] = 32'hFFFFFFF1;
    // rom_array[42922] = 32'hFFFFFFF1;
    // rom_array[42923] = 32'hFFFFFFF1;
    // rom_array[42924] = 32'hFFFFFFF1;
    // rom_array[42925] = 32'hFFFFFFF0;
    // rom_array[42926] = 32'hFFFFFFF0;
    // rom_array[42927] = 32'hFFFFFFF0;
    // rom_array[42928] = 32'hFFFFFFF0;
    // rom_array[42929] = 32'hFFFFFFF1;
    // rom_array[42930] = 32'hFFFFFFF1;
    // rom_array[42931] = 32'hFFFFFFF1;
    // rom_array[42932] = 32'hFFFFFFF1;
    // rom_array[42933] = 32'hFFFFFFF0;
    // rom_array[42934] = 32'hFFFFFFF0;
    // rom_array[42935] = 32'hFFFFFFF0;
    // rom_array[42936] = 32'hFFFFFFF0;
    // rom_array[42937] = 32'hFFFFFFF1;
    // rom_array[42938] = 32'hFFFFFFF1;
    // rom_array[42939] = 32'hFFFFFFF1;
    // rom_array[42940] = 32'hFFFFFFF1;
    // rom_array[42941] = 32'hFFFFFFF0;
    // rom_array[42942] = 32'hFFFFFFF0;
    // rom_array[42943] = 32'hFFFFFFF0;
    // rom_array[42944] = 32'hFFFFFFF0;
    // rom_array[42945] = 32'hFFFFFFF1;
    // rom_array[42946] = 32'hFFFFFFF1;
    // rom_array[42947] = 32'hFFFFFFF1;
    // rom_array[42948] = 32'hFFFFFFF1;
    // rom_array[42949] = 32'hFFFFFFF0;
    // rom_array[42950] = 32'hFFFFFFF0;
    // rom_array[42951] = 32'hFFFFFFF0;
    // rom_array[42952] = 32'hFFFFFFF0;
    // rom_array[42953] = 32'hFFFFFFF1;
    // rom_array[42954] = 32'hFFFFFFF1;
    // rom_array[42955] = 32'hFFFFFFF1;
    // rom_array[42956] = 32'hFFFFFFF1;
    // rom_array[42957] = 32'hFFFFFFF0;
    // rom_array[42958] = 32'hFFFFFFF0;
    // rom_array[42959] = 32'hFFFFFFF0;
    // rom_array[42960] = 32'hFFFFFFF0;
    // rom_array[42961] = 32'hFFFFFFF1;
    // rom_array[42962] = 32'hFFFFFFF1;
    // rom_array[42963] = 32'hFFFFFFF1;
    // rom_array[42964] = 32'hFFFFFFF1;
    // rom_array[42965] = 32'hFFFFFFF0;
    // rom_array[42966] = 32'hFFFFFFF0;
    // rom_array[42967] = 32'hFFFFFFF0;
    // rom_array[42968] = 32'hFFFFFFF0;
    // rom_array[42969] = 32'hFFFFFFF1;
    // rom_array[42970] = 32'hFFFFFFF1;
    // rom_array[42971] = 32'hFFFFFFF1;
    // rom_array[42972] = 32'hFFFFFFF1;
    // rom_array[42973] = 32'hFFFFFFF0;
    // rom_array[42974] = 32'hFFFFFFF0;
    // rom_array[42975] = 32'hFFFFFFF1;
    // rom_array[42976] = 32'hFFFFFFF1;
    // rom_array[42977] = 32'hFFFFFFF1;
    // rom_array[42978] = 32'hFFFFFFF1;
    // rom_array[42979] = 32'hFFFFFFF1;
    // rom_array[42980] = 32'hFFFFFFF1;
    // rom_array[42981] = 32'hFFFFFFF0;
    // rom_array[42982] = 32'hFFFFFFF0;
    // rom_array[42983] = 32'hFFFFFFF1;
    // rom_array[42984] = 32'hFFFFFFF1;
    // rom_array[42985] = 32'hFFFFFFF1;
    // rom_array[42986] = 32'hFFFFFFF1;
    // rom_array[42987] = 32'hFFFFFFF1;
    // rom_array[42988] = 32'hFFFFFFF1;
    // rom_array[42989] = 32'hFFFFFFF1;
    // rom_array[42990] = 32'hFFFFFFF1;
    // rom_array[42991] = 32'hFFFFFFF1;
    // rom_array[42992] = 32'hFFFFFFF1;
    // rom_array[42993] = 32'hFFFFFFF1;
    // rom_array[42994] = 32'hFFFFFFF1;
    // rom_array[42995] = 32'hFFFFFFF1;
    // rom_array[42996] = 32'hFFFFFFF1;
    // rom_array[42997] = 32'hFFFFFFF1;
    // rom_array[42998] = 32'hFFFFFFF1;
    // rom_array[42999] = 32'hFFFFFFF1;
    // rom_array[43000] = 32'hFFFFFFF1;
    // rom_array[43001] = 32'hFFFFFFF0;
    // rom_array[43002] = 32'hFFFFFFF0;
    // rom_array[43003] = 32'hFFFFFFF1;
    // rom_array[43004] = 32'hFFFFFFF1;
    // rom_array[43005] = 32'hFFFFFFF0;
    // rom_array[43006] = 32'hFFFFFFF0;
    // rom_array[43007] = 32'hFFFFFFF1;
    // rom_array[43008] = 32'hFFFFFFF1;
    // rom_array[43009] = 32'hFFFFFFF0;
    // rom_array[43010] = 32'hFFFFFFF0;
    // rom_array[43011] = 32'hFFFFFFF1;
    // rom_array[43012] = 32'hFFFFFFF1;
    // rom_array[43013] = 32'hFFFFFFF0;
    // rom_array[43014] = 32'hFFFFFFF0;
    // rom_array[43015] = 32'hFFFFFFF1;
    // rom_array[43016] = 32'hFFFFFFF1;
    // rom_array[43017] = 32'hFFFFFFF0;
    // rom_array[43018] = 32'hFFFFFFF0;
    // rom_array[43019] = 32'hFFFFFFF0;
    // rom_array[43020] = 32'hFFFFFFF0;
    // rom_array[43021] = 32'hFFFFFFF1;
    // rom_array[43022] = 32'hFFFFFFF1;
    // rom_array[43023] = 32'hFFFFFFF1;
    // rom_array[43024] = 32'hFFFFFFF1;
    // rom_array[43025] = 32'hFFFFFFF0;
    // rom_array[43026] = 32'hFFFFFFF0;
    // rom_array[43027] = 32'hFFFFFFF0;
    // rom_array[43028] = 32'hFFFFFFF0;
    // rom_array[43029] = 32'hFFFFFFF1;
    // rom_array[43030] = 32'hFFFFFFF1;
    // rom_array[43031] = 32'hFFFFFFF1;
    // rom_array[43032] = 32'hFFFFFFF1;
    // rom_array[43033] = 32'hFFFFFFF0;
    // rom_array[43034] = 32'hFFFFFFF0;
    // rom_array[43035] = 32'hFFFFFFF0;
    // rom_array[43036] = 32'hFFFFFFF0;
    // rom_array[43037] = 32'hFFFFFFF1;
    // rom_array[43038] = 32'hFFFFFFF1;
    // rom_array[43039] = 32'hFFFFFFF1;
    // rom_array[43040] = 32'hFFFFFFF1;
    // rom_array[43041] = 32'hFFFFFFF0;
    // rom_array[43042] = 32'hFFFFFFF0;
    // rom_array[43043] = 32'hFFFFFFF0;
    // rom_array[43044] = 32'hFFFFFFF0;
    // rom_array[43045] = 32'hFFFFFFF1;
    // rom_array[43046] = 32'hFFFFFFF1;
    // rom_array[43047] = 32'hFFFFFFF1;
    // rom_array[43048] = 32'hFFFFFFF1;
    // rom_array[43049] = 32'hFFFFFFF0;
    // rom_array[43050] = 32'hFFFFFFF0;
    // rom_array[43051] = 32'hFFFFFFF0;
    // rom_array[43052] = 32'hFFFFFFF0;
    // rom_array[43053] = 32'hFFFFFFF1;
    // rom_array[43054] = 32'hFFFFFFF1;
    // rom_array[43055] = 32'hFFFFFFF1;
    // rom_array[43056] = 32'hFFFFFFF1;
    // rom_array[43057] = 32'hFFFFFFF0;
    // rom_array[43058] = 32'hFFFFFFF0;
    // rom_array[43059] = 32'hFFFFFFF0;
    // rom_array[43060] = 32'hFFFFFFF0;
    // rom_array[43061] = 32'hFFFFFFF1;
    // rom_array[43062] = 32'hFFFFFFF1;
    // rom_array[43063] = 32'hFFFFFFF1;
    // rom_array[43064] = 32'hFFFFFFF1;
    // rom_array[43065] = 32'hFFFFFFF1;
    // rom_array[43066] = 32'hFFFFFFF1;
    // rom_array[43067] = 32'hFFFFFFF1;
    // rom_array[43068] = 32'hFFFFFFF1;
    // rom_array[43069] = 32'hFFFFFFF1;
    // rom_array[43070] = 32'hFFFFFFF1;
    // rom_array[43071] = 32'hFFFFFFF1;
    // rom_array[43072] = 32'hFFFFFFF1;
    // rom_array[43073] = 32'hFFFFFFF1;
    // rom_array[43074] = 32'hFFFFFFF1;
    // rom_array[43075] = 32'hFFFFFFF1;
    // rom_array[43076] = 32'hFFFFFFF1;
    // rom_array[43077] = 32'hFFFFFFF1;
    // rom_array[43078] = 32'hFFFFFFF1;
    // rom_array[43079] = 32'hFFFFFFF1;
    // rom_array[43080] = 32'hFFFFFFF1;
    // rom_array[43081] = 32'hFFFFFFF1;
    // rom_array[43082] = 32'hFFFFFFF1;
    // rom_array[43083] = 32'hFFFFFFF1;
    // rom_array[43084] = 32'hFFFFFFF1;
    // rom_array[43085] = 32'hFFFFFFF1;
    // rom_array[43086] = 32'hFFFFFFF1;
    // rom_array[43087] = 32'hFFFFFFF1;
    // rom_array[43088] = 32'hFFFFFFF1;
    // rom_array[43089] = 32'hFFFFFFF1;
    // rom_array[43090] = 32'hFFFFFFF1;
    // rom_array[43091] = 32'hFFFFFFF1;
    // rom_array[43092] = 32'hFFFFFFF1;
    // rom_array[43093] = 32'hFFFFFFF1;
    // rom_array[43094] = 32'hFFFFFFF1;
    // rom_array[43095] = 32'hFFFFFFF1;
    // rom_array[43096] = 32'hFFFFFFF1;
    // rom_array[43097] = 32'hFFFFFFF1;
    // rom_array[43098] = 32'hFFFFFFF1;
    // rom_array[43099] = 32'hFFFFFFF1;
    // rom_array[43100] = 32'hFFFFFFF1;
    // rom_array[43101] = 32'hFFFFFFF1;
    // rom_array[43102] = 32'hFFFFFFF1;
    // rom_array[43103] = 32'hFFFFFFF1;
    // rom_array[43104] = 32'hFFFFFFF1;
    // rom_array[43105] = 32'hFFFFFFF1;
    // rom_array[43106] = 32'hFFFFFFF1;
    // rom_array[43107] = 32'hFFFFFFF1;
    // rom_array[43108] = 32'hFFFFFFF1;
    // rom_array[43109] = 32'hFFFFFFF1;
    // rom_array[43110] = 32'hFFFFFFF1;
    // rom_array[43111] = 32'hFFFFFFF1;
    // rom_array[43112] = 32'hFFFFFFF1;
    // rom_array[43113] = 32'hFFFFFFF1;
    // rom_array[43114] = 32'hFFFFFFF1;
    // rom_array[43115] = 32'hFFFFFFF1;
    // rom_array[43116] = 32'hFFFFFFF1;
    // rom_array[43117] = 32'hFFFFFFF1;
    // rom_array[43118] = 32'hFFFFFFF1;
    // rom_array[43119] = 32'hFFFFFFF1;
    // rom_array[43120] = 32'hFFFFFFF1;
    // rom_array[43121] = 32'hFFFFFFF1;
    // rom_array[43122] = 32'hFFFFFFF1;
    // rom_array[43123] = 32'hFFFFFFF1;
    // rom_array[43124] = 32'hFFFFFFF1;
    // rom_array[43125] = 32'hFFFFFFF1;
    // rom_array[43126] = 32'hFFFFFFF1;
    // rom_array[43127] = 32'hFFFFFFF1;
    // rom_array[43128] = 32'hFFFFFFF1;
    // rom_array[43129] = 32'hFFFFFFF1;
    // rom_array[43130] = 32'hFFFFFFF1;
    // rom_array[43131] = 32'hFFFFFFF1;
    // rom_array[43132] = 32'hFFFFFFF1;
    // rom_array[43133] = 32'hFFFFFFF1;
    // rom_array[43134] = 32'hFFFFFFF1;
    // rom_array[43135] = 32'hFFFFFFF1;
    // rom_array[43136] = 32'hFFFFFFF1;
    // rom_array[43137] = 32'hFFFFFFF1;
    // rom_array[43138] = 32'hFFFFFFF1;
    // rom_array[43139] = 32'hFFFFFFF1;
    // rom_array[43140] = 32'hFFFFFFF1;
    // rom_array[43141] = 32'hFFFFFFF1;
    // rom_array[43142] = 32'hFFFFFFF1;
    // rom_array[43143] = 32'hFFFFFFF1;
    // rom_array[43144] = 32'hFFFFFFF1;
    // rom_array[43145] = 32'hFFFFFFF1;
    // rom_array[43146] = 32'hFFFFFFF1;
    // rom_array[43147] = 32'hFFFFFFF1;
    // rom_array[43148] = 32'hFFFFFFF1;
    // rom_array[43149] = 32'hFFFFFFF1;
    // rom_array[43150] = 32'hFFFFFFF1;
    // rom_array[43151] = 32'hFFFFFFF1;
    // rom_array[43152] = 32'hFFFFFFF1;
    // rom_array[43153] = 32'hFFFFFFF1;
    // rom_array[43154] = 32'hFFFFFFF1;
    // rom_array[43155] = 32'hFFFFFFF1;
    // rom_array[43156] = 32'hFFFFFFF1;
    // rom_array[43157] = 32'hFFFFFFF1;
    // rom_array[43158] = 32'hFFFFFFF1;
    // rom_array[43159] = 32'hFFFFFFF1;
    // rom_array[43160] = 32'hFFFFFFF1;
    // rom_array[43161] = 32'hFFFFFFF1;
    // rom_array[43162] = 32'hFFFFFFF1;
    // rom_array[43163] = 32'hFFFFFFF1;
    // rom_array[43164] = 32'hFFFFFFF1;
    // rom_array[43165] = 32'hFFFFFFF1;
    // rom_array[43166] = 32'hFFFFFFF1;
    // rom_array[43167] = 32'hFFFFFFF1;
    // rom_array[43168] = 32'hFFFFFFF1;
    // rom_array[43169] = 32'hFFFFFFF1;
    // rom_array[43170] = 32'hFFFFFFF1;
    // rom_array[43171] = 32'hFFFFFFF1;
    // rom_array[43172] = 32'hFFFFFFF1;
    // rom_array[43173] = 32'hFFFFFFF1;
    // rom_array[43174] = 32'hFFFFFFF1;
    // rom_array[43175] = 32'hFFFFFFF1;
    // rom_array[43176] = 32'hFFFFFFF1;
    // rom_array[43177] = 32'hFFFFFFF1;
    // rom_array[43178] = 32'hFFFFFFF1;
    // rom_array[43179] = 32'hFFFFFFF1;
    // rom_array[43180] = 32'hFFFFFFF1;
    // rom_array[43181] = 32'hFFFFFFF1;
    // rom_array[43182] = 32'hFFFFFFF1;
    // rom_array[43183] = 32'hFFFFFFF1;
    // rom_array[43184] = 32'hFFFFFFF1;
    // rom_array[43185] = 32'hFFFFFFF1;
    // rom_array[43186] = 32'hFFFFFFF1;
    // rom_array[43187] = 32'hFFFFFFF1;
    // rom_array[43188] = 32'hFFFFFFF1;
    // rom_array[43189] = 32'hFFFFFFF1;
    // rom_array[43190] = 32'hFFFFFFF1;
    // rom_array[43191] = 32'hFFFFFFF1;
    // rom_array[43192] = 32'hFFFFFFF1;
    // rom_array[43193] = 32'hFFFFFFF1;
    // rom_array[43194] = 32'hFFFFFFF1;
    // rom_array[43195] = 32'hFFFFFFF1;
    // rom_array[43196] = 32'hFFFFFFF1;
    // rom_array[43197] = 32'hFFFFFFF1;
    // rom_array[43198] = 32'hFFFFFFF1;
    // rom_array[43199] = 32'hFFFFFFF1;
    // rom_array[43200] = 32'hFFFFFFF1;
    // rom_array[43201] = 32'hFFFFFFF1;
    // rom_array[43202] = 32'hFFFFFFF1;
    // rom_array[43203] = 32'hFFFFFFF1;
    // rom_array[43204] = 32'hFFFFFFF1;
    // rom_array[43205] = 32'hFFFFFFF1;
    // rom_array[43206] = 32'hFFFFFFF1;
    // rom_array[43207] = 32'hFFFFFFF1;
    // rom_array[43208] = 32'hFFFFFFF1;
    // rom_array[43209] = 32'hFFFFFFF1;
    // rom_array[43210] = 32'hFFFFFFF1;
    // rom_array[43211] = 32'hFFFFFFF1;
    // rom_array[43212] = 32'hFFFFFFF1;
    // rom_array[43213] = 32'hFFFFFFF1;
    // rom_array[43214] = 32'hFFFFFFF1;
    // rom_array[43215] = 32'hFFFFFFF1;
    // rom_array[43216] = 32'hFFFFFFF1;
    // rom_array[43217] = 32'hFFFFFFF1;
    // rom_array[43218] = 32'hFFFFFFF1;
    // rom_array[43219] = 32'hFFFFFFF1;
    // rom_array[43220] = 32'hFFFFFFF1;
    // rom_array[43221] = 32'hFFFFFFF1;
    // rom_array[43222] = 32'hFFFFFFF1;
    // rom_array[43223] = 32'hFFFFFFF1;
    // rom_array[43224] = 32'hFFFFFFF1;
    // rom_array[43225] = 32'hFFFFFFF1;
    // rom_array[43226] = 32'hFFFFFFF1;
    // rom_array[43227] = 32'hFFFFFFF1;
    // rom_array[43228] = 32'hFFFFFFF1;
    // rom_array[43229] = 32'hFFFFFFF1;
    // rom_array[43230] = 32'hFFFFFFF1;
    // rom_array[43231] = 32'hFFFFFFF1;
    // rom_array[43232] = 32'hFFFFFFF1;
    // rom_array[43233] = 32'hFFFFFFF1;
    // rom_array[43234] = 32'hFFFFFFF1;
    // rom_array[43235] = 32'hFFFFFFF1;
    // rom_array[43236] = 32'hFFFFFFF1;
    // rom_array[43237] = 32'hFFFFFFF1;
    // rom_array[43238] = 32'hFFFFFFF1;
    // rom_array[43239] = 32'hFFFFFFF1;
    // rom_array[43240] = 32'hFFFFFFF1;
    // rom_array[43241] = 32'hFFFFFFF0;
    // rom_array[43242] = 32'hFFFFFFF0;
    // rom_array[43243] = 32'hFFFFFFF1;
    // rom_array[43244] = 32'hFFFFFFF1;
    // rom_array[43245] = 32'hFFFFFFF0;
    // rom_array[43246] = 32'hFFFFFFF0;
    // rom_array[43247] = 32'hFFFFFFF1;
    // rom_array[43248] = 32'hFFFFFFF1;
    // rom_array[43249] = 32'hFFFFFFF0;
    // rom_array[43250] = 32'hFFFFFFF0;
    // rom_array[43251] = 32'hFFFFFFF1;
    // rom_array[43252] = 32'hFFFFFFF1;
    // rom_array[43253] = 32'hFFFFFFF0;
    // rom_array[43254] = 32'hFFFFFFF0;
    // rom_array[43255] = 32'hFFFFFFF1;
    // rom_array[43256] = 32'hFFFFFFF1;
    // rom_array[43257] = 32'hFFFFFFF0;
    // rom_array[43258] = 32'hFFFFFFF0;
    // rom_array[43259] = 32'hFFFFFFF1;
    // rom_array[43260] = 32'hFFFFFFF1;
    // rom_array[43261] = 32'hFFFFFFF0;
    // rom_array[43262] = 32'hFFFFFFF0;
    // rom_array[43263] = 32'hFFFFFFF1;
    // rom_array[43264] = 32'hFFFFFFF1;
    // rom_array[43265] = 32'hFFFFFFF0;
    // rom_array[43266] = 32'hFFFFFFF0;
    // rom_array[43267] = 32'hFFFFFFF1;
    // rom_array[43268] = 32'hFFFFFFF1;
    // rom_array[43269] = 32'hFFFFFFF0;
    // rom_array[43270] = 32'hFFFFFFF0;
    // rom_array[43271] = 32'hFFFFFFF1;
    // rom_array[43272] = 32'hFFFFFFF1;
    // rom_array[43273] = 32'hFFFFFFF0;
    // rom_array[43274] = 32'hFFFFFFF0;
    // rom_array[43275] = 32'hFFFFFFF1;
    // rom_array[43276] = 32'hFFFFFFF1;
    // rom_array[43277] = 32'hFFFFFFF0;
    // rom_array[43278] = 32'hFFFFFFF0;
    // rom_array[43279] = 32'hFFFFFFF1;
    // rom_array[43280] = 32'hFFFFFFF1;
    // rom_array[43281] = 32'hFFFFFFF0;
    // rom_array[43282] = 32'hFFFFFFF0;
    // rom_array[43283] = 32'hFFFFFFF1;
    // rom_array[43284] = 32'hFFFFFFF1;
    // rom_array[43285] = 32'hFFFFFFF0;
    // rom_array[43286] = 32'hFFFFFFF0;
    // rom_array[43287] = 32'hFFFFFFF1;
    // rom_array[43288] = 32'hFFFFFFF1;
    // rom_array[43289] = 32'hFFFFFFF0;
    // rom_array[43290] = 32'hFFFFFFF0;
    // rom_array[43291] = 32'hFFFFFFF1;
    // rom_array[43292] = 32'hFFFFFFF1;
    // rom_array[43293] = 32'hFFFFFFF0;
    // rom_array[43294] = 32'hFFFFFFF0;
    // rom_array[43295] = 32'hFFFFFFF1;
    // rom_array[43296] = 32'hFFFFFFF1;
    // rom_array[43297] = 32'hFFFFFFF0;
    // rom_array[43298] = 32'hFFFFFFF0;
    // rom_array[43299] = 32'hFFFFFFF1;
    // rom_array[43300] = 32'hFFFFFFF1;
    // rom_array[43301] = 32'hFFFFFFF0;
    // rom_array[43302] = 32'hFFFFFFF0;
    // rom_array[43303] = 32'hFFFFFFF1;
    // rom_array[43304] = 32'hFFFFFFF1;
    // rom_array[43305] = 32'hFFFFFFF1;
    // rom_array[43306] = 32'hFFFFFFF1;
    // rom_array[43307] = 32'hFFFFFFF1;
    // rom_array[43308] = 32'hFFFFFFF1;
    // rom_array[43309] = 32'hFFFFFFF1;
    // rom_array[43310] = 32'hFFFFFFF1;
    // rom_array[43311] = 32'hFFFFFFF1;
    // rom_array[43312] = 32'hFFFFFFF1;
    // rom_array[43313] = 32'hFFFFFFF1;
    // rom_array[43314] = 32'hFFFFFFF1;
    // rom_array[43315] = 32'hFFFFFFF1;
    // rom_array[43316] = 32'hFFFFFFF1;
    // rom_array[43317] = 32'hFFFFFFF1;
    // rom_array[43318] = 32'hFFFFFFF1;
    // rom_array[43319] = 32'hFFFFFFF1;
    // rom_array[43320] = 32'hFFFFFFF1;
    // rom_array[43321] = 32'hFFFFFFF1;
    // rom_array[43322] = 32'hFFFFFFF1;
    // rom_array[43323] = 32'hFFFFFFF1;
    // rom_array[43324] = 32'hFFFFFFF1;
    // rom_array[43325] = 32'hFFFFFFF1;
    // rom_array[43326] = 32'hFFFFFFF1;
    // rom_array[43327] = 32'hFFFFFFF1;
    // rom_array[43328] = 32'hFFFFFFF1;
    // rom_array[43329] = 32'hFFFFFFF1;
    // rom_array[43330] = 32'hFFFFFFF1;
    // rom_array[43331] = 32'hFFFFFFF1;
    // rom_array[43332] = 32'hFFFFFFF1;
    // rom_array[43333] = 32'hFFFFFFF1;
    // rom_array[43334] = 32'hFFFFFFF1;
    // rom_array[43335] = 32'hFFFFFFF1;
    // rom_array[43336] = 32'hFFFFFFF1;
    // rom_array[43337] = 32'hFFFFFFF0;
    // rom_array[43338] = 32'hFFFFFFF0;
    // rom_array[43339] = 32'hFFFFFFF0;
    // rom_array[43340] = 32'hFFFFFFF0;
    // rom_array[43341] = 32'hFFFFFFF1;
    // rom_array[43342] = 32'hFFFFFFF1;
    // rom_array[43343] = 32'hFFFFFFF1;
    // rom_array[43344] = 32'hFFFFFFF1;
    // rom_array[43345] = 32'hFFFFFFF0;
    // rom_array[43346] = 32'hFFFFFFF0;
    // rom_array[43347] = 32'hFFFFFFF0;
    // rom_array[43348] = 32'hFFFFFFF0;
    // rom_array[43349] = 32'hFFFFFFF1;
    // rom_array[43350] = 32'hFFFFFFF1;
    // rom_array[43351] = 32'hFFFFFFF1;
    // rom_array[43352] = 32'hFFFFFFF1;
    // rom_array[43353] = 32'hFFFFFFF0;
    // rom_array[43354] = 32'hFFFFFFF0;
    // rom_array[43355] = 32'hFFFFFFF0;
    // rom_array[43356] = 32'hFFFFFFF0;
    // rom_array[43357] = 32'hFFFFFFF1;
    // rom_array[43358] = 32'hFFFFFFF1;
    // rom_array[43359] = 32'hFFFFFFF1;
    // rom_array[43360] = 32'hFFFFFFF1;
    // rom_array[43361] = 32'hFFFFFFF0;
    // rom_array[43362] = 32'hFFFFFFF0;
    // rom_array[43363] = 32'hFFFFFFF0;
    // rom_array[43364] = 32'hFFFFFFF0;
    // rom_array[43365] = 32'hFFFFFFF1;
    // rom_array[43366] = 32'hFFFFFFF1;
    // rom_array[43367] = 32'hFFFFFFF1;
    // rom_array[43368] = 32'hFFFFFFF1;
    // rom_array[43369] = 32'hFFFFFFF0;
    // rom_array[43370] = 32'hFFFFFFF0;
    // rom_array[43371] = 32'hFFFFFFF0;
    // rom_array[43372] = 32'hFFFFFFF0;
    // rom_array[43373] = 32'hFFFFFFF1;
    // rom_array[43374] = 32'hFFFFFFF1;
    // rom_array[43375] = 32'hFFFFFFF1;
    // rom_array[43376] = 32'hFFFFFFF1;
    // rom_array[43377] = 32'hFFFFFFF0;
    // rom_array[43378] = 32'hFFFFFFF0;
    // rom_array[43379] = 32'hFFFFFFF0;
    // rom_array[43380] = 32'hFFFFFFF0;
    // rom_array[43381] = 32'hFFFFFFF1;
    // rom_array[43382] = 32'hFFFFFFF1;
    // rom_array[43383] = 32'hFFFFFFF1;
    // rom_array[43384] = 32'hFFFFFFF1;
    // rom_array[43385] = 32'hFFFFFFF1;
    // rom_array[43386] = 32'hFFFFFFF1;
    // rom_array[43387] = 32'hFFFFFFF1;
    // rom_array[43388] = 32'hFFFFFFF1;
    // rom_array[43389] = 32'hFFFFFFF0;
    // rom_array[43390] = 32'hFFFFFFF0;
    // rom_array[43391] = 32'hFFFFFFF0;
    // rom_array[43392] = 32'hFFFFFFF0;
    // rom_array[43393] = 32'hFFFFFFF1;
    // rom_array[43394] = 32'hFFFFFFF1;
    // rom_array[43395] = 32'hFFFFFFF1;
    // rom_array[43396] = 32'hFFFFFFF1;
    // rom_array[43397] = 32'hFFFFFFF0;
    // rom_array[43398] = 32'hFFFFFFF0;
    // rom_array[43399] = 32'hFFFFFFF0;
    // rom_array[43400] = 32'hFFFFFFF0;
    // rom_array[43401] = 32'hFFFFFFF0;
    // rom_array[43402] = 32'hFFFFFFF0;
    // rom_array[43403] = 32'hFFFFFFF0;
    // rom_array[43404] = 32'hFFFFFFF0;
    // rom_array[43405] = 32'hFFFFFFF1;
    // rom_array[43406] = 32'hFFFFFFF1;
    // rom_array[43407] = 32'hFFFFFFF1;
    // rom_array[43408] = 32'hFFFFFFF1;
    // rom_array[43409] = 32'hFFFFFFF0;
    // rom_array[43410] = 32'hFFFFFFF0;
    // rom_array[43411] = 32'hFFFFFFF0;
    // rom_array[43412] = 32'hFFFFFFF0;
    // rom_array[43413] = 32'hFFFFFFF1;
    // rom_array[43414] = 32'hFFFFFFF1;
    // rom_array[43415] = 32'hFFFFFFF1;
    // rom_array[43416] = 32'hFFFFFFF1;
    // rom_array[43417] = 32'hFFFFFFF0;
    // rom_array[43418] = 32'hFFFFFFF0;
    // rom_array[43419] = 32'hFFFFFFF0;
    // rom_array[43420] = 32'hFFFFFFF0;
    // rom_array[43421] = 32'hFFFFFFF1;
    // rom_array[43422] = 32'hFFFFFFF1;
    // rom_array[43423] = 32'hFFFFFFF1;
    // rom_array[43424] = 32'hFFFFFFF1;
    // rom_array[43425] = 32'hFFFFFFF0;
    // rom_array[43426] = 32'hFFFFFFF0;
    // rom_array[43427] = 32'hFFFFFFF0;
    // rom_array[43428] = 32'hFFFFFFF0;
    // rom_array[43429] = 32'hFFFFFFF1;
    // rom_array[43430] = 32'hFFFFFFF1;
    // rom_array[43431] = 32'hFFFFFFF1;
    // rom_array[43432] = 32'hFFFFFFF1;
    // rom_array[43433] = 32'hFFFFFFF0;
    // rom_array[43434] = 32'hFFFFFFF0;
    // rom_array[43435] = 32'hFFFFFFF1;
    // rom_array[43436] = 32'hFFFFFFF1;
    // rom_array[43437] = 32'hFFFFFFF0;
    // rom_array[43438] = 32'hFFFFFFF0;
    // rom_array[43439] = 32'hFFFFFFF1;
    // rom_array[43440] = 32'hFFFFFFF1;
    // rom_array[43441] = 32'hFFFFFFF0;
    // rom_array[43442] = 32'hFFFFFFF0;
    // rom_array[43443] = 32'hFFFFFFF1;
    // rom_array[43444] = 32'hFFFFFFF1;
    // rom_array[43445] = 32'hFFFFFFF0;
    // rom_array[43446] = 32'hFFFFFFF0;
    // rom_array[43447] = 32'hFFFFFFF1;
    // rom_array[43448] = 32'hFFFFFFF1;
    // rom_array[43449] = 32'hFFFFFFF0;
    // rom_array[43450] = 32'hFFFFFFF0;
    // rom_array[43451] = 32'hFFFFFFF1;
    // rom_array[43452] = 32'hFFFFFFF1;
    // rom_array[43453] = 32'hFFFFFFF1;
    // rom_array[43454] = 32'hFFFFFFF1;
    // rom_array[43455] = 32'hFFFFFFF1;
    // rom_array[43456] = 32'hFFFFFFF1;
    // rom_array[43457] = 32'hFFFFFFF0;
    // rom_array[43458] = 32'hFFFFFFF0;
    // rom_array[43459] = 32'hFFFFFFF1;
    // rom_array[43460] = 32'hFFFFFFF1;
    // rom_array[43461] = 32'hFFFFFFF1;
    // rom_array[43462] = 32'hFFFFFFF1;
    // rom_array[43463] = 32'hFFFFFFF1;
    // rom_array[43464] = 32'hFFFFFFF1;
    // rom_array[43465] = 32'hFFFFFFF0;
    // rom_array[43466] = 32'hFFFFFFF0;
    // rom_array[43467] = 32'hFFFFFFF0;
    // rom_array[43468] = 32'hFFFFFFF0;
    // rom_array[43469] = 32'hFFFFFFF1;
    // rom_array[43470] = 32'hFFFFFFF1;
    // rom_array[43471] = 32'hFFFFFFF1;
    // rom_array[43472] = 32'hFFFFFFF1;
    // rom_array[43473] = 32'hFFFFFFF0;
    // rom_array[43474] = 32'hFFFFFFF0;
    // rom_array[43475] = 32'hFFFFFFF0;
    // rom_array[43476] = 32'hFFFFFFF0;
    // rom_array[43477] = 32'hFFFFFFF1;
    // rom_array[43478] = 32'hFFFFFFF1;
    // rom_array[43479] = 32'hFFFFFFF1;
    // rom_array[43480] = 32'hFFFFFFF1;
    // rom_array[43481] = 32'hFFFFFFF0;
    // rom_array[43482] = 32'hFFFFFFF0;
    // rom_array[43483] = 32'hFFFFFFF1;
    // rom_array[43484] = 32'hFFFFFFF1;
    // rom_array[43485] = 32'hFFFFFFF0;
    // rom_array[43486] = 32'hFFFFFFF0;
    // rom_array[43487] = 32'hFFFFFFF0;
    // rom_array[43488] = 32'hFFFFFFF0;
    // rom_array[43489] = 32'hFFFFFFF0;
    // rom_array[43490] = 32'hFFFFFFF0;
    // rom_array[43491] = 32'hFFFFFFF1;
    // rom_array[43492] = 32'hFFFFFFF1;
    // rom_array[43493] = 32'hFFFFFFF0;
    // rom_array[43494] = 32'hFFFFFFF0;
    // rom_array[43495] = 32'hFFFFFFF0;
    // rom_array[43496] = 32'hFFFFFFF0;
    // rom_array[43497] = 32'hFFFFFFF1;
    // rom_array[43498] = 32'hFFFFFFF1;
    // rom_array[43499] = 32'hFFFFFFF1;
    // rom_array[43500] = 32'hFFFFFFF1;
    // rom_array[43501] = 32'hFFFFFFF1;
    // rom_array[43502] = 32'hFFFFFFF1;
    // rom_array[43503] = 32'hFFFFFFF1;
    // rom_array[43504] = 32'hFFFFFFF1;
    // rom_array[43505] = 32'hFFFFFFF1;
    // rom_array[43506] = 32'hFFFFFFF1;
    // rom_array[43507] = 32'hFFFFFFF1;
    // rom_array[43508] = 32'hFFFFFFF1;
    // rom_array[43509] = 32'hFFFFFFF1;
    // rom_array[43510] = 32'hFFFFFFF1;
    // rom_array[43511] = 32'hFFFFFFF1;
    // rom_array[43512] = 32'hFFFFFFF1;
    // rom_array[43513] = 32'hFFFFFFF1;
    // rom_array[43514] = 32'hFFFFFFF1;
    // rom_array[43515] = 32'hFFFFFFF1;
    // rom_array[43516] = 32'hFFFFFFF1;
    // rom_array[43517] = 32'hFFFFFFF1;
    // rom_array[43518] = 32'hFFFFFFF1;
    // rom_array[43519] = 32'hFFFFFFF1;
    // rom_array[43520] = 32'hFFFFFFF1;
    // rom_array[43521] = 32'hFFFFFFF1;
    // rom_array[43522] = 32'hFFFFFFF1;
    // rom_array[43523] = 32'hFFFFFFF1;
    // rom_array[43524] = 32'hFFFFFFF1;
    // rom_array[43525] = 32'hFFFFFFF1;
    // rom_array[43526] = 32'hFFFFFFF1;
    // rom_array[43527] = 32'hFFFFFFF1;
    // rom_array[43528] = 32'hFFFFFFF1;
    // rom_array[43529] = 32'hFFFFFFF1;
    // rom_array[43530] = 32'hFFFFFFF1;
    // rom_array[43531] = 32'hFFFFFFF1;
    // rom_array[43532] = 32'hFFFFFFF1;
    // rom_array[43533] = 32'hFFFFFFF1;
    // rom_array[43534] = 32'hFFFFFFF1;
    // rom_array[43535] = 32'hFFFFFFF1;
    // rom_array[43536] = 32'hFFFFFFF1;
    // rom_array[43537] = 32'hFFFFFFF1;
    // rom_array[43538] = 32'hFFFFFFF1;
    // rom_array[43539] = 32'hFFFFFFF1;
    // rom_array[43540] = 32'hFFFFFFF1;
    // rom_array[43541] = 32'hFFFFFFF1;
    // rom_array[43542] = 32'hFFFFFFF1;
    // rom_array[43543] = 32'hFFFFFFF1;
    // rom_array[43544] = 32'hFFFFFFF1;
    // rom_array[43545] = 32'hFFFFFFF1;
    // rom_array[43546] = 32'hFFFFFFF1;
    // rom_array[43547] = 32'hFFFFFFF1;
    // rom_array[43548] = 32'hFFFFFFF1;
    // rom_array[43549] = 32'hFFFFFFF1;
    // rom_array[43550] = 32'hFFFFFFF1;
    // rom_array[43551] = 32'hFFFFFFF1;
    // rom_array[43552] = 32'hFFFFFFF1;
    // rom_array[43553] = 32'hFFFFFFF1;
    // rom_array[43554] = 32'hFFFFFFF1;
    // rom_array[43555] = 32'hFFFFFFF1;
    // rom_array[43556] = 32'hFFFFFFF1;
    // rom_array[43557] = 32'hFFFFFFF1;
    // rom_array[43558] = 32'hFFFFFFF1;
    // rom_array[43559] = 32'hFFFFFFF1;
    // rom_array[43560] = 32'hFFFFFFF1;
    // rom_array[43561] = 32'hFFFFFFF1;
    // rom_array[43562] = 32'hFFFFFFF1;
    // rom_array[43563] = 32'hFFFFFFF1;
    // rom_array[43564] = 32'hFFFFFFF1;
    // rom_array[43565] = 32'hFFFFFFF1;
    // rom_array[43566] = 32'hFFFFFFF1;
    // rom_array[43567] = 32'hFFFFFFF1;
    // rom_array[43568] = 32'hFFFFFFF1;
    // rom_array[43569] = 32'hFFFFFFF1;
    // rom_array[43570] = 32'hFFFFFFF1;
    // rom_array[43571] = 32'hFFFFFFF1;
    // rom_array[43572] = 32'hFFFFFFF1;
    // rom_array[43573] = 32'hFFFFFFF1;
    // rom_array[43574] = 32'hFFFFFFF1;
    // rom_array[43575] = 32'hFFFFFFF1;
    // rom_array[43576] = 32'hFFFFFFF1;
    // rom_array[43577] = 32'hFFFFFFF1;
    // rom_array[43578] = 32'hFFFFFFF1;
    // rom_array[43579] = 32'hFFFFFFF1;
    // rom_array[43580] = 32'hFFFFFFF1;
    // rom_array[43581] = 32'hFFFFFFF1;
    // rom_array[43582] = 32'hFFFFFFF1;
    // rom_array[43583] = 32'hFFFFFFF1;
    // rom_array[43584] = 32'hFFFFFFF1;
    // rom_array[43585] = 32'hFFFFFFF1;
    // rom_array[43586] = 32'hFFFFFFF1;
    // rom_array[43587] = 32'hFFFFFFF1;
    // rom_array[43588] = 32'hFFFFFFF1;
    // rom_array[43589] = 32'hFFFFFFF1;
    // rom_array[43590] = 32'hFFFFFFF1;
    // rom_array[43591] = 32'hFFFFFFF1;
    // rom_array[43592] = 32'hFFFFFFF1;
    // rom_array[43593] = 32'hFFFFFFF1;
    // rom_array[43594] = 32'hFFFFFFF1;
    // rom_array[43595] = 32'hFFFFFFF1;
    // rom_array[43596] = 32'hFFFFFFF1;
    // rom_array[43597] = 32'hFFFFFFF1;
    // rom_array[43598] = 32'hFFFFFFF1;
    // rom_array[43599] = 32'hFFFFFFF1;
    // rom_array[43600] = 32'hFFFFFFF1;
    // rom_array[43601] = 32'hFFFFFFF1;
    // rom_array[43602] = 32'hFFFFFFF1;
    // rom_array[43603] = 32'hFFFFFFF1;
    // rom_array[43604] = 32'hFFFFFFF1;
    // rom_array[43605] = 32'hFFFFFFF1;
    // rom_array[43606] = 32'hFFFFFFF1;
    // rom_array[43607] = 32'hFFFFFFF1;
    // rom_array[43608] = 32'hFFFFFFF1;
    // rom_array[43609] = 32'hFFFFFFF1;
    // rom_array[43610] = 32'hFFFFFFF1;
    // rom_array[43611] = 32'hFFFFFFF1;
    // rom_array[43612] = 32'hFFFFFFF1;
    // rom_array[43613] = 32'hFFFFFFF1;
    // rom_array[43614] = 32'hFFFFFFF1;
    // rom_array[43615] = 32'hFFFFFFF1;
    // rom_array[43616] = 32'hFFFFFFF1;
    // rom_array[43617] = 32'hFFFFFFF1;
    // rom_array[43618] = 32'hFFFFFFF1;
    // rom_array[43619] = 32'hFFFFFFF1;
    // rom_array[43620] = 32'hFFFFFFF1;
    // rom_array[43621] = 32'hFFFFFFF1;
    // rom_array[43622] = 32'hFFFFFFF1;
    // rom_array[43623] = 32'hFFFFFFF1;
    // rom_array[43624] = 32'hFFFFFFF1;
    // rom_array[43625] = 32'hFFFFFFF1;
    // rom_array[43626] = 32'hFFFFFFF1;
    // rom_array[43627] = 32'hFFFFFFF1;
    // rom_array[43628] = 32'hFFFFFFF1;
    // rom_array[43629] = 32'hFFFFFFF0;
    // rom_array[43630] = 32'hFFFFFFF0;
    // rom_array[43631] = 32'hFFFFFFF0;
    // rom_array[43632] = 32'hFFFFFFF0;
    // rom_array[43633] = 32'hFFFFFFF1;
    // rom_array[43634] = 32'hFFFFFFF1;
    // rom_array[43635] = 32'hFFFFFFF1;
    // rom_array[43636] = 32'hFFFFFFF1;
    // rom_array[43637] = 32'hFFFFFFF0;
    // rom_array[43638] = 32'hFFFFFFF0;
    // rom_array[43639] = 32'hFFFFFFF0;
    // rom_array[43640] = 32'hFFFFFFF0;
    // rom_array[43641] = 32'hFFFFFFF1;
    // rom_array[43642] = 32'hFFFFFFF1;
    // rom_array[43643] = 32'hFFFFFFF1;
    // rom_array[43644] = 32'hFFFFFFF1;
    // rom_array[43645] = 32'hFFFFFFF0;
    // rom_array[43646] = 32'hFFFFFFF0;
    // rom_array[43647] = 32'hFFFFFFF0;
    // rom_array[43648] = 32'hFFFFFFF0;
    // rom_array[43649] = 32'hFFFFFFF1;
    // rom_array[43650] = 32'hFFFFFFF1;
    // rom_array[43651] = 32'hFFFFFFF1;
    // rom_array[43652] = 32'hFFFFFFF1;
    // rom_array[43653] = 32'hFFFFFFF0;
    // rom_array[43654] = 32'hFFFFFFF0;
    // rom_array[43655] = 32'hFFFFFFF0;
    // rom_array[43656] = 32'hFFFFFFF0;
    // rom_array[43657] = 32'hFFFFFFF1;
    // rom_array[43658] = 32'hFFFFFFF1;
    // rom_array[43659] = 32'hFFFFFFF1;
    // rom_array[43660] = 32'hFFFFFFF1;
    // rom_array[43661] = 32'hFFFFFFF0;
    // rom_array[43662] = 32'hFFFFFFF0;
    // rom_array[43663] = 32'hFFFFFFF0;
    // rom_array[43664] = 32'hFFFFFFF0;
    // rom_array[43665] = 32'hFFFFFFF1;
    // rom_array[43666] = 32'hFFFFFFF1;
    // rom_array[43667] = 32'hFFFFFFF1;
    // rom_array[43668] = 32'hFFFFFFF1;
    // rom_array[43669] = 32'hFFFFFFF0;
    // rom_array[43670] = 32'hFFFFFFF0;
    // rom_array[43671] = 32'hFFFFFFF0;
    // rom_array[43672] = 32'hFFFFFFF0;
    // rom_array[43673] = 32'hFFFFFFF1;
    // rom_array[43674] = 32'hFFFFFFF1;
    // rom_array[43675] = 32'hFFFFFFF1;
    // rom_array[43676] = 32'hFFFFFFF1;
    // rom_array[43677] = 32'hFFFFFFF0;
    // rom_array[43678] = 32'hFFFFFFF0;
    // rom_array[43679] = 32'hFFFFFFF0;
    // rom_array[43680] = 32'hFFFFFFF0;
    // rom_array[43681] = 32'hFFFFFFF1;
    // rom_array[43682] = 32'hFFFFFFF1;
    // rom_array[43683] = 32'hFFFFFFF1;
    // rom_array[43684] = 32'hFFFFFFF1;
    // rom_array[43685] = 32'hFFFFFFF0;
    // rom_array[43686] = 32'hFFFFFFF0;
    // rom_array[43687] = 32'hFFFFFFF0;
    // rom_array[43688] = 32'hFFFFFFF0;
    // rom_array[43689] = 32'hFFFFFFF1;
    // rom_array[43690] = 32'hFFFFFFF1;
    // rom_array[43691] = 32'hFFFFFFF1;
    // rom_array[43692] = 32'hFFFFFFF1;
    // rom_array[43693] = 32'hFFFFFFF0;
    // rom_array[43694] = 32'hFFFFFFF0;
    // rom_array[43695] = 32'hFFFFFFF0;
    // rom_array[43696] = 32'hFFFFFFF0;
    // rom_array[43697] = 32'hFFFFFFF1;
    // rom_array[43698] = 32'hFFFFFFF1;
    // rom_array[43699] = 32'hFFFFFFF1;
    // rom_array[43700] = 32'hFFFFFFF1;
    // rom_array[43701] = 32'hFFFFFFF0;
    // rom_array[43702] = 32'hFFFFFFF0;
    // rom_array[43703] = 32'hFFFFFFF0;
    // rom_array[43704] = 32'hFFFFFFF0;
    // rom_array[43705] = 32'hFFFFFFF1;
    // rom_array[43706] = 32'hFFFFFFF1;
    // rom_array[43707] = 32'hFFFFFFF1;
    // rom_array[43708] = 32'hFFFFFFF1;
    // rom_array[43709] = 32'hFFFFFFF0;
    // rom_array[43710] = 32'hFFFFFFF0;
    // rom_array[43711] = 32'hFFFFFFF0;
    // rom_array[43712] = 32'hFFFFFFF0;
    // rom_array[43713] = 32'hFFFFFFF1;
    // rom_array[43714] = 32'hFFFFFFF1;
    // rom_array[43715] = 32'hFFFFFFF1;
    // rom_array[43716] = 32'hFFFFFFF1;
    // rom_array[43717] = 32'hFFFFFFF0;
    // rom_array[43718] = 32'hFFFFFFF0;
    // rom_array[43719] = 32'hFFFFFFF0;
    // rom_array[43720] = 32'hFFFFFFF0;
    // rom_array[43721] = 32'hFFFFFFF1;
    // rom_array[43722] = 32'hFFFFFFF1;
    // rom_array[43723] = 32'hFFFFFFF1;
    // rom_array[43724] = 32'hFFFFFFF1;
    // rom_array[43725] = 32'hFFFFFFF0;
    // rom_array[43726] = 32'hFFFFFFF0;
    // rom_array[43727] = 32'hFFFFFFF0;
    // rom_array[43728] = 32'hFFFFFFF0;
    // rom_array[43729] = 32'hFFFFFFF1;
    // rom_array[43730] = 32'hFFFFFFF1;
    // rom_array[43731] = 32'hFFFFFFF1;
    // rom_array[43732] = 32'hFFFFFFF1;
    // rom_array[43733] = 32'hFFFFFFF0;
    // rom_array[43734] = 32'hFFFFFFF0;
    // rom_array[43735] = 32'hFFFFFFF0;
    // rom_array[43736] = 32'hFFFFFFF0;
    // rom_array[43737] = 32'hFFFFFFF1;
    // rom_array[43738] = 32'hFFFFFFF1;
    // rom_array[43739] = 32'hFFFFFFF1;
    // rom_array[43740] = 32'hFFFFFFF1;
    // rom_array[43741] = 32'hFFFFFFF0;
    // rom_array[43742] = 32'hFFFFFFF0;
    // rom_array[43743] = 32'hFFFFFFF0;
    // rom_array[43744] = 32'hFFFFFFF0;
    // rom_array[43745] = 32'hFFFFFFF1;
    // rom_array[43746] = 32'hFFFFFFF1;
    // rom_array[43747] = 32'hFFFFFFF1;
    // rom_array[43748] = 32'hFFFFFFF1;
    // rom_array[43749] = 32'hFFFFFFF0;
    // rom_array[43750] = 32'hFFFFFFF0;
    // rom_array[43751] = 32'hFFFFFFF0;
    // rom_array[43752] = 32'hFFFFFFF0;
    // rom_array[43753] = 32'hFFFFFFF1;
    // rom_array[43754] = 32'hFFFFFFF1;
    // rom_array[43755] = 32'hFFFFFFF1;
    // rom_array[43756] = 32'hFFFFFFF1;
    // rom_array[43757] = 32'hFFFFFFF0;
    // rom_array[43758] = 32'hFFFFFFF0;
    // rom_array[43759] = 32'hFFFFFFF0;
    // rom_array[43760] = 32'hFFFFFFF0;
    // rom_array[43761] = 32'hFFFFFFF1;
    // rom_array[43762] = 32'hFFFFFFF1;
    // rom_array[43763] = 32'hFFFFFFF1;
    // rom_array[43764] = 32'hFFFFFFF1;
    // rom_array[43765] = 32'hFFFFFFF0;
    // rom_array[43766] = 32'hFFFFFFF0;
    // rom_array[43767] = 32'hFFFFFFF0;
    // rom_array[43768] = 32'hFFFFFFF0;
    // rom_array[43769] = 32'hFFFFFFF1;
    // rom_array[43770] = 32'hFFFFFFF1;
    // rom_array[43771] = 32'hFFFFFFF1;
    // rom_array[43772] = 32'hFFFFFFF1;
    // rom_array[43773] = 32'hFFFFFFF1;
    // rom_array[43774] = 32'hFFFFFFF1;
    // rom_array[43775] = 32'hFFFFFFF1;
    // rom_array[43776] = 32'hFFFFFFF1;
    // rom_array[43777] = 32'hFFFFFFF1;
    // rom_array[43778] = 32'hFFFFFFF1;
    // rom_array[43779] = 32'hFFFFFFF1;
    // rom_array[43780] = 32'hFFFFFFF1;
    // rom_array[43781] = 32'hFFFFFFF1;
    // rom_array[43782] = 32'hFFFFFFF1;
    // rom_array[43783] = 32'hFFFFFFF1;
    // rom_array[43784] = 32'hFFFFFFF1;
    // rom_array[43785] = 32'hFFFFFFF1;
    // rom_array[43786] = 32'hFFFFFFF1;
    // rom_array[43787] = 32'hFFFFFFF1;
    // rom_array[43788] = 32'hFFFFFFF1;
    // rom_array[43789] = 32'hFFFFFFF0;
    // rom_array[43790] = 32'hFFFFFFF0;
    // rom_array[43791] = 32'hFFFFFFF0;
    // rom_array[43792] = 32'hFFFFFFF0;
    // rom_array[43793] = 32'hFFFFFFF1;
    // rom_array[43794] = 32'hFFFFFFF1;
    // rom_array[43795] = 32'hFFFFFFF1;
    // rom_array[43796] = 32'hFFFFFFF1;
    // rom_array[43797] = 32'hFFFFFFF0;
    // rom_array[43798] = 32'hFFFFFFF0;
    // rom_array[43799] = 32'hFFFFFFF0;
    // rom_array[43800] = 32'hFFFFFFF0;
    // rom_array[43801] = 32'hFFFFFFF1;
    // rom_array[43802] = 32'hFFFFFFF1;
    // rom_array[43803] = 32'hFFFFFFF1;
    // rom_array[43804] = 32'hFFFFFFF1;
    // rom_array[43805] = 32'hFFFFFFF0;
    // rom_array[43806] = 32'hFFFFFFF0;
    // rom_array[43807] = 32'hFFFFFFF0;
    // rom_array[43808] = 32'hFFFFFFF0;
    // rom_array[43809] = 32'hFFFFFFF1;
    // rom_array[43810] = 32'hFFFFFFF1;
    // rom_array[43811] = 32'hFFFFFFF1;
    // rom_array[43812] = 32'hFFFFFFF1;
    // rom_array[43813] = 32'hFFFFFFF0;
    // rom_array[43814] = 32'hFFFFFFF0;
    // rom_array[43815] = 32'hFFFFFFF0;
    // rom_array[43816] = 32'hFFFFFFF0;
    // rom_array[43817] = 32'hFFFFFFF0;
    // rom_array[43818] = 32'hFFFFFFF0;
    // rom_array[43819] = 32'hFFFFFFF0;
    // rom_array[43820] = 32'hFFFFFFF0;
    // rom_array[43821] = 32'hFFFFFFF0;
    // rom_array[43822] = 32'hFFFFFFF0;
    // rom_array[43823] = 32'hFFFFFFF1;
    // rom_array[43824] = 32'hFFFFFFF1;
    // rom_array[43825] = 32'hFFFFFFF0;
    // rom_array[43826] = 32'hFFFFFFF0;
    // rom_array[43827] = 32'hFFFFFFF0;
    // rom_array[43828] = 32'hFFFFFFF0;
    // rom_array[43829] = 32'hFFFFFFF0;
    // rom_array[43830] = 32'hFFFFFFF0;
    // rom_array[43831] = 32'hFFFFFFF1;
    // rom_array[43832] = 32'hFFFFFFF1;
    // rom_array[43833] = 32'hFFFFFFF0;
    // rom_array[43834] = 32'hFFFFFFF0;
    // rom_array[43835] = 32'hFFFFFFF0;
    // rom_array[43836] = 32'hFFFFFFF0;
    // rom_array[43837] = 32'hFFFFFFF1;
    // rom_array[43838] = 32'hFFFFFFF1;
    // rom_array[43839] = 32'hFFFFFFF1;
    // rom_array[43840] = 32'hFFFFFFF1;
    // rom_array[43841] = 32'hFFFFFFF0;
    // rom_array[43842] = 32'hFFFFFFF0;
    // rom_array[43843] = 32'hFFFFFFF0;
    // rom_array[43844] = 32'hFFFFFFF0;
    // rom_array[43845] = 32'hFFFFFFF1;
    // rom_array[43846] = 32'hFFFFFFF1;
    // rom_array[43847] = 32'hFFFFFFF1;
    // rom_array[43848] = 32'hFFFFFFF1;
    // rom_array[43849] = 32'hFFFFFFF0;
    // rom_array[43850] = 32'hFFFFFFF0;
    // rom_array[43851] = 32'hFFFFFFF1;
    // rom_array[43852] = 32'hFFFFFFF1;
    // rom_array[43853] = 32'hFFFFFFF0;
    // rom_array[43854] = 32'hFFFFFFF0;
    // rom_array[43855] = 32'hFFFFFFF1;
    // rom_array[43856] = 32'hFFFFFFF1;
    // rom_array[43857] = 32'hFFFFFFF0;
    // rom_array[43858] = 32'hFFFFFFF0;
    // rom_array[43859] = 32'hFFFFFFF1;
    // rom_array[43860] = 32'hFFFFFFF1;
    // rom_array[43861] = 32'hFFFFFFF0;
    // rom_array[43862] = 32'hFFFFFFF0;
    // rom_array[43863] = 32'hFFFFFFF1;
    // rom_array[43864] = 32'hFFFFFFF1;
    // rom_array[43865] = 32'hFFFFFFF0;
    // rom_array[43866] = 32'hFFFFFFF0;
    // rom_array[43867] = 32'hFFFFFFF1;
    // rom_array[43868] = 32'hFFFFFFF1;
    // rom_array[43869] = 32'hFFFFFFF0;
    // rom_array[43870] = 32'hFFFFFFF0;
    // rom_array[43871] = 32'hFFFFFFF1;
    // rom_array[43872] = 32'hFFFFFFF1;
    // rom_array[43873] = 32'hFFFFFFF0;
    // rom_array[43874] = 32'hFFFFFFF0;
    // rom_array[43875] = 32'hFFFFFFF1;
    // rom_array[43876] = 32'hFFFFFFF1;
    // rom_array[43877] = 32'hFFFFFFF0;
    // rom_array[43878] = 32'hFFFFFFF0;
    // rom_array[43879] = 32'hFFFFFFF1;
    // rom_array[43880] = 32'hFFFFFFF1;
    // rom_array[43881] = 32'hFFFFFFF0;
    // rom_array[43882] = 32'hFFFFFFF0;
    // rom_array[43883] = 32'hFFFFFFF0;
    // rom_array[43884] = 32'hFFFFFFF0;
    // rom_array[43885] = 32'hFFFFFFF1;
    // rom_array[43886] = 32'hFFFFFFF1;
    // rom_array[43887] = 32'hFFFFFFF1;
    // rom_array[43888] = 32'hFFFFFFF1;
    // rom_array[43889] = 32'hFFFFFFF0;
    // rom_array[43890] = 32'hFFFFFFF0;
    // rom_array[43891] = 32'hFFFFFFF0;
    // rom_array[43892] = 32'hFFFFFFF0;
    // rom_array[43893] = 32'hFFFFFFF1;
    // rom_array[43894] = 32'hFFFFFFF1;
    // rom_array[43895] = 32'hFFFFFFF1;
    // rom_array[43896] = 32'hFFFFFFF1;
    // rom_array[43897] = 32'hFFFFFFF0;
    // rom_array[43898] = 32'hFFFFFFF0;
    // rom_array[43899] = 32'hFFFFFFF0;
    // rom_array[43900] = 32'hFFFFFFF0;
    // rom_array[43901] = 32'hFFFFFFF1;
    // rom_array[43902] = 32'hFFFFFFF1;
    // rom_array[43903] = 32'hFFFFFFF1;
    // rom_array[43904] = 32'hFFFFFFF1;
    // rom_array[43905] = 32'hFFFFFFF0;
    // rom_array[43906] = 32'hFFFFFFF0;
    // rom_array[43907] = 32'hFFFFFFF0;
    // rom_array[43908] = 32'hFFFFFFF0;
    // rom_array[43909] = 32'hFFFFFFF1;
    // rom_array[43910] = 32'hFFFFFFF1;
    // rom_array[43911] = 32'hFFFFFFF1;
    // rom_array[43912] = 32'hFFFFFFF1;
    // rom_array[43913] = 32'hFFFFFFF0;
    // rom_array[43914] = 32'hFFFFFFF0;
    // rom_array[43915] = 32'hFFFFFFF0;
    // rom_array[43916] = 32'hFFFFFFF0;
    // rom_array[43917] = 32'hFFFFFFF1;
    // rom_array[43918] = 32'hFFFFFFF1;
    // rom_array[43919] = 32'hFFFFFFF1;
    // rom_array[43920] = 32'hFFFFFFF1;
    // rom_array[43921] = 32'hFFFFFFF0;
    // rom_array[43922] = 32'hFFFFFFF0;
    // rom_array[43923] = 32'hFFFFFFF0;
    // rom_array[43924] = 32'hFFFFFFF0;
    // rom_array[43925] = 32'hFFFFFFF1;
    // rom_array[43926] = 32'hFFFFFFF1;
    // rom_array[43927] = 32'hFFFFFFF1;
    // rom_array[43928] = 32'hFFFFFFF1;
    // rom_array[43929] = 32'hFFFFFFF0;
    // rom_array[43930] = 32'hFFFFFFF0;
    // rom_array[43931] = 32'hFFFFFFF0;
    // rom_array[43932] = 32'hFFFFFFF0;
    // rom_array[43933] = 32'hFFFFFFF1;
    // rom_array[43934] = 32'hFFFFFFF1;
    // rom_array[43935] = 32'hFFFFFFF1;
    // rom_array[43936] = 32'hFFFFFFF1;
    // rom_array[43937] = 32'hFFFFFFF0;
    // rom_array[43938] = 32'hFFFFFFF0;
    // rom_array[43939] = 32'hFFFFFFF0;
    // rom_array[43940] = 32'hFFFFFFF0;
    // rom_array[43941] = 32'hFFFFFFF1;
    // rom_array[43942] = 32'hFFFFFFF1;
    // rom_array[43943] = 32'hFFFFFFF1;
    // rom_array[43944] = 32'hFFFFFFF1;
    // rom_array[43945] = 32'hFFFFFFF0;
    // rom_array[43946] = 32'hFFFFFFF0;
    // rom_array[43947] = 32'hFFFFFFF1;
    // rom_array[43948] = 32'hFFFFFFF1;
    // rom_array[43949] = 32'hFFFFFFF0;
    // rom_array[43950] = 32'hFFFFFFF0;
    // rom_array[43951] = 32'hFFFFFFF1;
    // rom_array[43952] = 32'hFFFFFFF1;
    // rom_array[43953] = 32'hFFFFFFF0;
    // rom_array[43954] = 32'hFFFFFFF0;
    // rom_array[43955] = 32'hFFFFFFF1;
    // rom_array[43956] = 32'hFFFFFFF1;
    // rom_array[43957] = 32'hFFFFFFF0;
    // rom_array[43958] = 32'hFFFFFFF0;
    // rom_array[43959] = 32'hFFFFFFF1;
    // rom_array[43960] = 32'hFFFFFFF1;
    // rom_array[43961] = 32'hFFFFFFF0;
    // rom_array[43962] = 32'hFFFFFFF0;
    // rom_array[43963] = 32'hFFFFFFF1;
    // rom_array[43964] = 32'hFFFFFFF1;
    // rom_array[43965] = 32'hFFFFFFF0;
    // rom_array[43966] = 32'hFFFFFFF0;
    // rom_array[43967] = 32'hFFFFFFF1;
    // rom_array[43968] = 32'hFFFFFFF1;
    // rom_array[43969] = 32'hFFFFFFF0;
    // rom_array[43970] = 32'hFFFFFFF0;
    // rom_array[43971] = 32'hFFFFFFF1;
    // rom_array[43972] = 32'hFFFFFFF1;
    // rom_array[43973] = 32'hFFFFFFF0;
    // rom_array[43974] = 32'hFFFFFFF0;
    // rom_array[43975] = 32'hFFFFFFF1;
    // rom_array[43976] = 32'hFFFFFFF1;
    // rom_array[43977] = 32'hFFFFFFF0;
    // rom_array[43978] = 32'hFFFFFFF0;
    // rom_array[43979] = 32'hFFFFFFF0;
    // rom_array[43980] = 32'hFFFFFFF0;
    // rom_array[43981] = 32'hFFFFFFF1;
    // rom_array[43982] = 32'hFFFFFFF1;
    // rom_array[43983] = 32'hFFFFFFF1;
    // rom_array[43984] = 32'hFFFFFFF1;
    // rom_array[43985] = 32'hFFFFFFF0;
    // rom_array[43986] = 32'hFFFFFFF0;
    // rom_array[43987] = 32'hFFFFFFF0;
    // rom_array[43988] = 32'hFFFFFFF0;
    // rom_array[43989] = 32'hFFFFFFF1;
    // rom_array[43990] = 32'hFFFFFFF1;
    // rom_array[43991] = 32'hFFFFFFF1;
    // rom_array[43992] = 32'hFFFFFFF1;
    // rom_array[43993] = 32'hFFFFFFF0;
    // rom_array[43994] = 32'hFFFFFFF0;
    // rom_array[43995] = 32'hFFFFFFF0;
    // rom_array[43996] = 32'hFFFFFFF0;
    // rom_array[43997] = 32'hFFFFFFF1;
    // rom_array[43998] = 32'hFFFFFFF1;
    // rom_array[43999] = 32'hFFFFFFF1;
    // rom_array[44000] = 32'hFFFFFFF1;
    // rom_array[44001] = 32'hFFFFFFF0;
    // rom_array[44002] = 32'hFFFFFFF0;
    // rom_array[44003] = 32'hFFFFFFF0;
    // rom_array[44004] = 32'hFFFFFFF0;
    // rom_array[44005] = 32'hFFFFFFF1;
    // rom_array[44006] = 32'hFFFFFFF1;
    // rom_array[44007] = 32'hFFFFFFF1;
    // rom_array[44008] = 32'hFFFFFFF1;
    // rom_array[44009] = 32'hFFFFFFF0;
    // rom_array[44010] = 32'hFFFFFFF0;
    // rom_array[44011] = 32'hFFFFFFF1;
    // rom_array[44012] = 32'hFFFFFFF1;
    // rom_array[44013] = 32'hFFFFFFF1;
    // rom_array[44014] = 32'hFFFFFFF1;
    // rom_array[44015] = 32'hFFFFFFF1;
    // rom_array[44016] = 32'hFFFFFFF1;
    // rom_array[44017] = 32'hFFFFFFF0;
    // rom_array[44018] = 32'hFFFFFFF0;
    // rom_array[44019] = 32'hFFFFFFF1;
    // rom_array[44020] = 32'hFFFFFFF1;
    // rom_array[44021] = 32'hFFFFFFF1;
    // rom_array[44022] = 32'hFFFFFFF1;
    // rom_array[44023] = 32'hFFFFFFF1;
    // rom_array[44024] = 32'hFFFFFFF1;
    // rom_array[44025] = 32'hFFFFFFF1;
    // rom_array[44026] = 32'hFFFFFFF1;
    // rom_array[44027] = 32'hFFFFFFF1;
    // rom_array[44028] = 32'hFFFFFFF1;
    // rom_array[44029] = 32'hFFFFFFF1;
    // rom_array[44030] = 32'hFFFFFFF1;
    // rom_array[44031] = 32'hFFFFFFF1;
    // rom_array[44032] = 32'hFFFFFFF1;
    // rom_array[44033] = 32'hFFFFFFF1;
    // rom_array[44034] = 32'hFFFFFFF1;
    // rom_array[44035] = 32'hFFFFFFF1;
    // rom_array[44036] = 32'hFFFFFFF1;
    // rom_array[44037] = 32'hFFFFFFF1;
    // rom_array[44038] = 32'hFFFFFFF1;
    // rom_array[44039] = 32'hFFFFFFF1;
    // rom_array[44040] = 32'hFFFFFFF1;
    // rom_array[44041] = 32'hFFFFFFF0;
    // rom_array[44042] = 32'hFFFFFFF0;
    // rom_array[44043] = 32'hFFFFFFF0;
    // rom_array[44044] = 32'hFFFFFFF0;
    // rom_array[44045] = 32'hFFFFFFF1;
    // rom_array[44046] = 32'hFFFFFFF1;
    // rom_array[44047] = 32'hFFFFFFF1;
    // rom_array[44048] = 32'hFFFFFFF1;
    // rom_array[44049] = 32'hFFFFFFF0;
    // rom_array[44050] = 32'hFFFFFFF0;
    // rom_array[44051] = 32'hFFFFFFF0;
    // rom_array[44052] = 32'hFFFFFFF0;
    // rom_array[44053] = 32'hFFFFFFF1;
    // rom_array[44054] = 32'hFFFFFFF1;
    // rom_array[44055] = 32'hFFFFFFF1;
    // rom_array[44056] = 32'hFFFFFFF1;
    // rom_array[44057] = 32'hFFFFFFF0;
    // rom_array[44058] = 32'hFFFFFFF0;
    // rom_array[44059] = 32'hFFFFFFF0;
    // rom_array[44060] = 32'hFFFFFFF0;
    // rom_array[44061] = 32'hFFFFFFF1;
    // rom_array[44062] = 32'hFFFFFFF1;
    // rom_array[44063] = 32'hFFFFFFF1;
    // rom_array[44064] = 32'hFFFFFFF1;
    // rom_array[44065] = 32'hFFFFFFF0;
    // rom_array[44066] = 32'hFFFFFFF0;
    // rom_array[44067] = 32'hFFFFFFF0;
    // rom_array[44068] = 32'hFFFFFFF0;
    // rom_array[44069] = 32'hFFFFFFF1;
    // rom_array[44070] = 32'hFFFFFFF1;
    // rom_array[44071] = 32'hFFFFFFF1;
    // rom_array[44072] = 32'hFFFFFFF1;
    // rom_array[44073] = 32'hFFFFFFF0;
    // rom_array[44074] = 32'hFFFFFFF0;
    // rom_array[44075] = 32'hFFFFFFF0;
    // rom_array[44076] = 32'hFFFFFFF0;
    // rom_array[44077] = 32'hFFFFFFF1;
    // rom_array[44078] = 32'hFFFFFFF1;
    // rom_array[44079] = 32'hFFFFFFF1;
    // rom_array[44080] = 32'hFFFFFFF1;
    // rom_array[44081] = 32'hFFFFFFF0;
    // rom_array[44082] = 32'hFFFFFFF0;
    // rom_array[44083] = 32'hFFFFFFF0;
    // rom_array[44084] = 32'hFFFFFFF0;
    // rom_array[44085] = 32'hFFFFFFF1;
    // rom_array[44086] = 32'hFFFFFFF1;
    // rom_array[44087] = 32'hFFFFFFF1;
    // rom_array[44088] = 32'hFFFFFFF1;
    // rom_array[44089] = 32'hFFFFFFF1;
    // rom_array[44090] = 32'hFFFFFFF1;
    // rom_array[44091] = 32'hFFFFFFF1;
    // rom_array[44092] = 32'hFFFFFFF1;
    // rom_array[44093] = 32'hFFFFFFF1;
    // rom_array[44094] = 32'hFFFFFFF1;
    // rom_array[44095] = 32'hFFFFFFF1;
    // rom_array[44096] = 32'hFFFFFFF1;
    // rom_array[44097] = 32'hFFFFFFF1;
    // rom_array[44098] = 32'hFFFFFFF1;
    // rom_array[44099] = 32'hFFFFFFF1;
    // rom_array[44100] = 32'hFFFFFFF1;
    // rom_array[44101] = 32'hFFFFFFF1;
    // rom_array[44102] = 32'hFFFFFFF1;
    // rom_array[44103] = 32'hFFFFFFF1;
    // rom_array[44104] = 32'hFFFFFFF1;
    // rom_array[44105] = 32'hFFFFFFF1;
    // rom_array[44106] = 32'hFFFFFFF1;
    // rom_array[44107] = 32'hFFFFFFF1;
    // rom_array[44108] = 32'hFFFFFFF1;
    // rom_array[44109] = 32'hFFFFFFF1;
    // rom_array[44110] = 32'hFFFFFFF1;
    // rom_array[44111] = 32'hFFFFFFF1;
    // rom_array[44112] = 32'hFFFFFFF1;
    // rom_array[44113] = 32'hFFFFFFF1;
    // rom_array[44114] = 32'hFFFFFFF1;
    // rom_array[44115] = 32'hFFFFFFF1;
    // rom_array[44116] = 32'hFFFFFFF1;
    // rom_array[44117] = 32'hFFFFFFF1;
    // rom_array[44118] = 32'hFFFFFFF1;
    // rom_array[44119] = 32'hFFFFFFF1;
    // rom_array[44120] = 32'hFFFFFFF1;
    // rom_array[44121] = 32'hFFFFFFF1;
    // rom_array[44122] = 32'hFFFFFFF1;
    // rom_array[44123] = 32'hFFFFFFF1;
    // rom_array[44124] = 32'hFFFFFFF1;
    // rom_array[44125] = 32'hFFFFFFF1;
    // rom_array[44126] = 32'hFFFFFFF1;
    // rom_array[44127] = 32'hFFFFFFF1;
    // rom_array[44128] = 32'hFFFFFFF1;
    // rom_array[44129] = 32'hFFFFFFF1;
    // rom_array[44130] = 32'hFFFFFFF1;
    // rom_array[44131] = 32'hFFFFFFF1;
    // rom_array[44132] = 32'hFFFFFFF1;
    // rom_array[44133] = 32'hFFFFFFF1;
    // rom_array[44134] = 32'hFFFFFFF1;
    // rom_array[44135] = 32'hFFFFFFF1;
    // rom_array[44136] = 32'hFFFFFFF1;
    // rom_array[44137] = 32'hFFFFFFF1;
    // rom_array[44138] = 32'hFFFFFFF1;
    // rom_array[44139] = 32'hFFFFFFF1;
    // rom_array[44140] = 32'hFFFFFFF1;
    // rom_array[44141] = 32'hFFFFFFF1;
    // rom_array[44142] = 32'hFFFFFFF1;
    // rom_array[44143] = 32'hFFFFFFF1;
    // rom_array[44144] = 32'hFFFFFFF1;
    // rom_array[44145] = 32'hFFFFFFF1;
    // rom_array[44146] = 32'hFFFFFFF1;
    // rom_array[44147] = 32'hFFFFFFF1;
    // rom_array[44148] = 32'hFFFFFFF1;
    // rom_array[44149] = 32'hFFFFFFF1;
    // rom_array[44150] = 32'hFFFFFFF1;
    // rom_array[44151] = 32'hFFFFFFF1;
    // rom_array[44152] = 32'hFFFFFFF1;
    // rom_array[44153] = 32'hFFFFFFF1;
    // rom_array[44154] = 32'hFFFFFFF1;
    // rom_array[44155] = 32'hFFFFFFF1;
    // rom_array[44156] = 32'hFFFFFFF1;
    // rom_array[44157] = 32'hFFFFFFF1;
    // rom_array[44158] = 32'hFFFFFFF1;
    // rom_array[44159] = 32'hFFFFFFF1;
    // rom_array[44160] = 32'hFFFFFFF1;
    // rom_array[44161] = 32'hFFFFFFF1;
    // rom_array[44162] = 32'hFFFFFFF1;
    // rom_array[44163] = 32'hFFFFFFF1;
    // rom_array[44164] = 32'hFFFFFFF1;
    // rom_array[44165] = 32'hFFFFFFF1;
    // rom_array[44166] = 32'hFFFFFFF1;
    // rom_array[44167] = 32'hFFFFFFF1;
    // rom_array[44168] = 32'hFFFFFFF1;
    // rom_array[44169] = 32'hFFFFFFF1;
    // rom_array[44170] = 32'hFFFFFFF1;
    // rom_array[44171] = 32'hFFFFFFF1;
    // rom_array[44172] = 32'hFFFFFFF1;
    // rom_array[44173] = 32'hFFFFFFF1;
    // rom_array[44174] = 32'hFFFFFFF1;
    // rom_array[44175] = 32'hFFFFFFF1;
    // rom_array[44176] = 32'hFFFFFFF1;
    // rom_array[44177] = 32'hFFFFFFF1;
    // rom_array[44178] = 32'hFFFFFFF1;
    // rom_array[44179] = 32'hFFFFFFF1;
    // rom_array[44180] = 32'hFFFFFFF1;
    // rom_array[44181] = 32'hFFFFFFF1;
    // rom_array[44182] = 32'hFFFFFFF1;
    // rom_array[44183] = 32'hFFFFFFF1;
    // rom_array[44184] = 32'hFFFFFFF1;
    // rom_array[44185] = 32'hFFFFFFF1;
    // rom_array[44186] = 32'hFFFFFFF1;
    // rom_array[44187] = 32'hFFFFFFF1;
    // rom_array[44188] = 32'hFFFFFFF1;
    // rom_array[44189] = 32'hFFFFFFF0;
    // rom_array[44190] = 32'hFFFFFFF0;
    // rom_array[44191] = 32'hFFFFFFF0;
    // rom_array[44192] = 32'hFFFFFFF0;
    // rom_array[44193] = 32'hFFFFFFF1;
    // rom_array[44194] = 32'hFFFFFFF1;
    // rom_array[44195] = 32'hFFFFFFF1;
    // rom_array[44196] = 32'hFFFFFFF1;
    // rom_array[44197] = 32'hFFFFFFF0;
    // rom_array[44198] = 32'hFFFFFFF0;
    // rom_array[44199] = 32'hFFFFFFF0;
    // rom_array[44200] = 32'hFFFFFFF0;
    // rom_array[44201] = 32'hFFFFFFF1;
    // rom_array[44202] = 32'hFFFFFFF1;
    // rom_array[44203] = 32'hFFFFFFF1;
    // rom_array[44204] = 32'hFFFFFFF1;
    // rom_array[44205] = 32'hFFFFFFF0;
    // rom_array[44206] = 32'hFFFFFFF0;
    // rom_array[44207] = 32'hFFFFFFF0;
    // rom_array[44208] = 32'hFFFFFFF0;
    // rom_array[44209] = 32'hFFFFFFF1;
    // rom_array[44210] = 32'hFFFFFFF1;
    // rom_array[44211] = 32'hFFFFFFF1;
    // rom_array[44212] = 32'hFFFFFFF1;
    // rom_array[44213] = 32'hFFFFFFF0;
    // rom_array[44214] = 32'hFFFFFFF0;
    // rom_array[44215] = 32'hFFFFFFF0;
    // rom_array[44216] = 32'hFFFFFFF0;
    // rom_array[44217] = 32'hFFFFFFF1;
    // rom_array[44218] = 32'hFFFFFFF1;
    // rom_array[44219] = 32'hFFFFFFF1;
    // rom_array[44220] = 32'hFFFFFFF1;
    // rom_array[44221] = 32'hFFFFFFF0;
    // rom_array[44222] = 32'hFFFFFFF0;
    // rom_array[44223] = 32'hFFFFFFF0;
    // rom_array[44224] = 32'hFFFFFFF0;
    // rom_array[44225] = 32'hFFFFFFF1;
    // rom_array[44226] = 32'hFFFFFFF1;
    // rom_array[44227] = 32'hFFFFFFF1;
    // rom_array[44228] = 32'hFFFFFFF1;
    // rom_array[44229] = 32'hFFFFFFF0;
    // rom_array[44230] = 32'hFFFFFFF0;
    // rom_array[44231] = 32'hFFFFFFF0;
    // rom_array[44232] = 32'hFFFFFFF0;
    // rom_array[44233] = 32'hFFFFFFF1;
    // rom_array[44234] = 32'hFFFFFFF1;
    // rom_array[44235] = 32'hFFFFFFF1;
    // rom_array[44236] = 32'hFFFFFFF1;
    // rom_array[44237] = 32'hFFFFFFF0;
    // rom_array[44238] = 32'hFFFFFFF0;
    // rom_array[44239] = 32'hFFFFFFF0;
    // rom_array[44240] = 32'hFFFFFFF0;
    // rom_array[44241] = 32'hFFFFFFF1;
    // rom_array[44242] = 32'hFFFFFFF1;
    // rom_array[44243] = 32'hFFFFFFF1;
    // rom_array[44244] = 32'hFFFFFFF1;
    // rom_array[44245] = 32'hFFFFFFF0;
    // rom_array[44246] = 32'hFFFFFFF0;
    // rom_array[44247] = 32'hFFFFFFF0;
    // rom_array[44248] = 32'hFFFFFFF0;
    // rom_array[44249] = 32'hFFFFFFF1;
    // rom_array[44250] = 32'hFFFFFFF1;
    // rom_array[44251] = 32'hFFFFFFF1;
    // rom_array[44252] = 32'hFFFFFFF1;
    // rom_array[44253] = 32'hFFFFFFF1;
    // rom_array[44254] = 32'hFFFFFFF1;
    // rom_array[44255] = 32'hFFFFFFF1;
    // rom_array[44256] = 32'hFFFFFFF1;
    // rom_array[44257] = 32'hFFFFFFF1;
    // rom_array[44258] = 32'hFFFFFFF1;
    // rom_array[44259] = 32'hFFFFFFF1;
    // rom_array[44260] = 32'hFFFFFFF1;
    // rom_array[44261] = 32'hFFFFFFF1;
    // rom_array[44262] = 32'hFFFFFFF1;
    // rom_array[44263] = 32'hFFFFFFF1;
    // rom_array[44264] = 32'hFFFFFFF1;
    // rom_array[44265] = 32'hFFFFFFF1;
    // rom_array[44266] = 32'hFFFFFFF1;
    // rom_array[44267] = 32'hFFFFFFF1;
    // rom_array[44268] = 32'hFFFFFFF1;
    // rom_array[44269] = 32'hFFFFFFF1;
    // rom_array[44270] = 32'hFFFFFFF1;
    // rom_array[44271] = 32'hFFFFFFF1;
    // rom_array[44272] = 32'hFFFFFFF1;
    // rom_array[44273] = 32'hFFFFFFF1;
    // rom_array[44274] = 32'hFFFFFFF1;
    // rom_array[44275] = 32'hFFFFFFF1;
    // rom_array[44276] = 32'hFFFFFFF1;
    // rom_array[44277] = 32'hFFFFFFF1;
    // rom_array[44278] = 32'hFFFFFFF1;
    // rom_array[44279] = 32'hFFFFFFF1;
    // rom_array[44280] = 32'hFFFFFFF1;
    // rom_array[44281] = 32'hFFFFFFF1;
    // rom_array[44282] = 32'hFFFFFFF1;
    // rom_array[44283] = 32'hFFFFFFF1;
    // rom_array[44284] = 32'hFFFFFFF1;
    // rom_array[44285] = 32'hFFFFFFF0;
    // rom_array[44286] = 32'hFFFFFFF0;
    // rom_array[44287] = 32'hFFFFFFF0;
    // rom_array[44288] = 32'hFFFFFFF0;
    // rom_array[44289] = 32'hFFFFFFF1;
    // rom_array[44290] = 32'hFFFFFFF1;
    // rom_array[44291] = 32'hFFFFFFF1;
    // rom_array[44292] = 32'hFFFFFFF1;
    // rom_array[44293] = 32'hFFFFFFF0;
    // rom_array[44294] = 32'hFFFFFFF0;
    // rom_array[44295] = 32'hFFFFFFF0;
    // rom_array[44296] = 32'hFFFFFFF0;
    // rom_array[44297] = 32'hFFFFFFF1;
    // rom_array[44298] = 32'hFFFFFFF1;
    // rom_array[44299] = 32'hFFFFFFF1;
    // rom_array[44300] = 32'hFFFFFFF1;
    // rom_array[44301] = 32'hFFFFFFF0;
    // rom_array[44302] = 32'hFFFFFFF0;
    // rom_array[44303] = 32'hFFFFFFF0;
    // rom_array[44304] = 32'hFFFFFFF0;
    // rom_array[44305] = 32'hFFFFFFF1;
    // rom_array[44306] = 32'hFFFFFFF1;
    // rom_array[44307] = 32'hFFFFFFF1;
    // rom_array[44308] = 32'hFFFFFFF1;
    // rom_array[44309] = 32'hFFFFFFF0;
    // rom_array[44310] = 32'hFFFFFFF0;
    // rom_array[44311] = 32'hFFFFFFF0;
    // rom_array[44312] = 32'hFFFFFFF0;
    // rom_array[44313] = 32'hFFFFFFF1;
    // rom_array[44314] = 32'hFFFFFFF1;
    // rom_array[44315] = 32'hFFFFFFF1;
    // rom_array[44316] = 32'hFFFFFFF1;
    // rom_array[44317] = 32'hFFFFFFF0;
    // rom_array[44318] = 32'hFFFFFFF0;
    // rom_array[44319] = 32'hFFFFFFF1;
    // rom_array[44320] = 32'hFFFFFFF1;
    // rom_array[44321] = 32'hFFFFFFF1;
    // rom_array[44322] = 32'hFFFFFFF1;
    // rom_array[44323] = 32'hFFFFFFF1;
    // rom_array[44324] = 32'hFFFFFFF1;
    // rom_array[44325] = 32'hFFFFFFF0;
    // rom_array[44326] = 32'hFFFFFFF0;
    // rom_array[44327] = 32'hFFFFFFF1;
    // rom_array[44328] = 32'hFFFFFFF1;
    // rom_array[44329] = 32'hFFFFFFF0;
    // rom_array[44330] = 32'hFFFFFFF0;
    // rom_array[44331] = 32'hFFFFFFF1;
    // rom_array[44332] = 32'hFFFFFFF1;
    // rom_array[44333] = 32'hFFFFFFF0;
    // rom_array[44334] = 32'hFFFFFFF0;
    // rom_array[44335] = 32'hFFFFFFF1;
    // rom_array[44336] = 32'hFFFFFFF1;
    // rom_array[44337] = 32'hFFFFFFF0;
    // rom_array[44338] = 32'hFFFFFFF0;
    // rom_array[44339] = 32'hFFFFFFF1;
    // rom_array[44340] = 32'hFFFFFFF1;
    // rom_array[44341] = 32'hFFFFFFF0;
    // rom_array[44342] = 32'hFFFFFFF0;
    // rom_array[44343] = 32'hFFFFFFF1;
    // rom_array[44344] = 32'hFFFFFFF1;
    // rom_array[44345] = 32'hFFFFFFF0;
    // rom_array[44346] = 32'hFFFFFFF0;
    // rom_array[44347] = 32'hFFFFFFF1;
    // rom_array[44348] = 32'hFFFFFFF1;
    // rom_array[44349] = 32'hFFFFFFF0;
    // rom_array[44350] = 32'hFFFFFFF0;
    // rom_array[44351] = 32'hFFFFFFF1;
    // rom_array[44352] = 32'hFFFFFFF1;
    // rom_array[44353] = 32'hFFFFFFF0;
    // rom_array[44354] = 32'hFFFFFFF0;
    // rom_array[44355] = 32'hFFFFFFF1;
    // rom_array[44356] = 32'hFFFFFFF1;
    // rom_array[44357] = 32'hFFFFFFF0;
    // rom_array[44358] = 32'hFFFFFFF0;
    // rom_array[44359] = 32'hFFFFFFF1;
    // rom_array[44360] = 32'hFFFFFFF1;
    // rom_array[44361] = 32'hFFFFFFF0;
    // rom_array[44362] = 32'hFFFFFFF0;
    // rom_array[44363] = 32'hFFFFFFF1;
    // rom_array[44364] = 32'hFFFFFFF1;
    // rom_array[44365] = 32'hFFFFFFF0;
    // rom_array[44366] = 32'hFFFFFFF0;
    // rom_array[44367] = 32'hFFFFFFF1;
    // rom_array[44368] = 32'hFFFFFFF1;
    // rom_array[44369] = 32'hFFFFFFF0;
    // rom_array[44370] = 32'hFFFFFFF0;
    // rom_array[44371] = 32'hFFFFFFF1;
    // rom_array[44372] = 32'hFFFFFFF1;
    // rom_array[44373] = 32'hFFFFFFF0;
    // rom_array[44374] = 32'hFFFFFFF0;
    // rom_array[44375] = 32'hFFFFFFF1;
    // rom_array[44376] = 32'hFFFFFFF1;
    // rom_array[44377] = 32'hFFFFFFF0;
    // rom_array[44378] = 32'hFFFFFFF0;
    // rom_array[44379] = 32'hFFFFFFF1;
    // rom_array[44380] = 32'hFFFFFFF1;
    // rom_array[44381] = 32'hFFFFFFF0;
    // rom_array[44382] = 32'hFFFFFFF0;
    // rom_array[44383] = 32'hFFFFFFF1;
    // rom_array[44384] = 32'hFFFFFFF1;
    // rom_array[44385] = 32'hFFFFFFF0;
    // rom_array[44386] = 32'hFFFFFFF0;
    // rom_array[44387] = 32'hFFFFFFF1;
    // rom_array[44388] = 32'hFFFFFFF1;
    // rom_array[44389] = 32'hFFFFFFF0;
    // rom_array[44390] = 32'hFFFFFFF0;
    // rom_array[44391] = 32'hFFFFFFF1;
    // rom_array[44392] = 32'hFFFFFFF1;
    // rom_array[44393] = 32'hFFFFFFF0;
    // rom_array[44394] = 32'hFFFFFFF0;
    // rom_array[44395] = 32'hFFFFFFF1;
    // rom_array[44396] = 32'hFFFFFFF1;
    // rom_array[44397] = 32'hFFFFFFF0;
    // rom_array[44398] = 32'hFFFFFFF0;
    // rom_array[44399] = 32'hFFFFFFF0;
    // rom_array[44400] = 32'hFFFFFFF0;
    // rom_array[44401] = 32'hFFFFFFF0;
    // rom_array[44402] = 32'hFFFFFFF0;
    // rom_array[44403] = 32'hFFFFFFF1;
    // rom_array[44404] = 32'hFFFFFFF1;
    // rom_array[44405] = 32'hFFFFFFF0;
    // rom_array[44406] = 32'hFFFFFFF0;
    // rom_array[44407] = 32'hFFFFFFF0;
    // rom_array[44408] = 32'hFFFFFFF0;
    // rom_array[44409] = 32'hFFFFFFF1;
    // rom_array[44410] = 32'hFFFFFFF1;
    // rom_array[44411] = 32'hFFFFFFF1;
    // rom_array[44412] = 32'hFFFFFFF1;
    // rom_array[44413] = 32'hFFFFFFF0;
    // rom_array[44414] = 32'hFFFFFFF0;
    // rom_array[44415] = 32'hFFFFFFF0;
    // rom_array[44416] = 32'hFFFFFFF0;
    // rom_array[44417] = 32'hFFFFFFF1;
    // rom_array[44418] = 32'hFFFFFFF1;
    // rom_array[44419] = 32'hFFFFFFF1;
    // rom_array[44420] = 32'hFFFFFFF1;
    // rom_array[44421] = 32'hFFFFFFF0;
    // rom_array[44422] = 32'hFFFFFFF0;
    // rom_array[44423] = 32'hFFFFFFF0;
    // rom_array[44424] = 32'hFFFFFFF0;
    // rom_array[44425] = 32'hFFFFFFF1;
    // rom_array[44426] = 32'hFFFFFFF1;
    // rom_array[44427] = 32'hFFFFFFF1;
    // rom_array[44428] = 32'hFFFFFFF1;
    // rom_array[44429] = 32'hFFFFFFF1;
    // rom_array[44430] = 32'hFFFFFFF1;
    // rom_array[44431] = 32'hFFFFFFF1;
    // rom_array[44432] = 32'hFFFFFFF1;
    // rom_array[44433] = 32'hFFFFFFF1;
    // rom_array[44434] = 32'hFFFFFFF1;
    // rom_array[44435] = 32'hFFFFFFF1;
    // rom_array[44436] = 32'hFFFFFFF1;
    // rom_array[44437] = 32'hFFFFFFF1;
    // rom_array[44438] = 32'hFFFFFFF1;
    // rom_array[44439] = 32'hFFFFFFF1;
    // rom_array[44440] = 32'hFFFFFFF1;
    // rom_array[44441] = 32'hFFFFFFF1;
    // rom_array[44442] = 32'hFFFFFFF1;
    // rom_array[44443] = 32'hFFFFFFF1;
    // rom_array[44444] = 32'hFFFFFFF1;
    // rom_array[44445] = 32'hFFFFFFF1;
    // rom_array[44446] = 32'hFFFFFFF1;
    // rom_array[44447] = 32'hFFFFFFF1;
    // rom_array[44448] = 32'hFFFFFFF1;
    // rom_array[44449] = 32'hFFFFFFF1;
    // rom_array[44450] = 32'hFFFFFFF1;
    // rom_array[44451] = 32'hFFFFFFF1;
    // rom_array[44452] = 32'hFFFFFFF1;
    // rom_array[44453] = 32'hFFFFFFF1;
    // rom_array[44454] = 32'hFFFFFFF1;
    // rom_array[44455] = 32'hFFFFFFF1;
    // rom_array[44456] = 32'hFFFFFFF1;
    // rom_array[44457] = 32'hFFFFFFF1;
    // rom_array[44458] = 32'hFFFFFFF1;
    // rom_array[44459] = 32'hFFFFFFF1;
    // rom_array[44460] = 32'hFFFFFFF1;
    // rom_array[44461] = 32'hFFFFFFF1;
    // rom_array[44462] = 32'hFFFFFFF1;
    // rom_array[44463] = 32'hFFFFFFF1;
    // rom_array[44464] = 32'hFFFFFFF1;
    // rom_array[44465] = 32'hFFFFFFF1;
    // rom_array[44466] = 32'hFFFFFFF1;
    // rom_array[44467] = 32'hFFFFFFF1;
    // rom_array[44468] = 32'hFFFFFFF1;
    // rom_array[44469] = 32'hFFFFFFF1;
    // rom_array[44470] = 32'hFFFFFFF1;
    // rom_array[44471] = 32'hFFFFFFF1;
    // rom_array[44472] = 32'hFFFFFFF1;
    // rom_array[44473] = 32'hFFFFFFF1;
    // rom_array[44474] = 32'hFFFFFFF1;
    // rom_array[44475] = 32'hFFFFFFF1;
    // rom_array[44476] = 32'hFFFFFFF1;
    // rom_array[44477] = 32'hFFFFFFF1;
    // rom_array[44478] = 32'hFFFFFFF1;
    // rom_array[44479] = 32'hFFFFFFF1;
    // rom_array[44480] = 32'hFFFFFFF1;
    // rom_array[44481] = 32'hFFFFFFF1;
    // rom_array[44482] = 32'hFFFFFFF1;
    // rom_array[44483] = 32'hFFFFFFF1;
    // rom_array[44484] = 32'hFFFFFFF1;
    // rom_array[44485] = 32'hFFFFFFF1;
    // rom_array[44486] = 32'hFFFFFFF1;
    // rom_array[44487] = 32'hFFFFFFF1;
    // rom_array[44488] = 32'hFFFFFFF1;
    // rom_array[44489] = 32'hFFFFFFF1;
    // rom_array[44490] = 32'hFFFFFFF1;
    // rom_array[44491] = 32'hFFFFFFF1;
    // rom_array[44492] = 32'hFFFFFFF1;
    // rom_array[44493] = 32'hFFFFFFF1;
    // rom_array[44494] = 32'hFFFFFFF1;
    // rom_array[44495] = 32'hFFFFFFF1;
    // rom_array[44496] = 32'hFFFFFFF1;
    // rom_array[44497] = 32'hFFFFFFF1;
    // rom_array[44498] = 32'hFFFFFFF1;
    // rom_array[44499] = 32'hFFFFFFF1;
    // rom_array[44500] = 32'hFFFFFFF1;
    // rom_array[44501] = 32'hFFFFFFF1;
    // rom_array[44502] = 32'hFFFFFFF1;
    // rom_array[44503] = 32'hFFFFFFF1;
    // rom_array[44504] = 32'hFFFFFFF1;
    // rom_array[44505] = 32'hFFFFFFF1;
    // rom_array[44506] = 32'hFFFFFFF1;
    // rom_array[44507] = 32'hFFFFFFF1;
    // rom_array[44508] = 32'hFFFFFFF1;
    // rom_array[44509] = 32'hFFFFFFF1;
    // rom_array[44510] = 32'hFFFFFFF1;
    // rom_array[44511] = 32'hFFFFFFF1;
    // rom_array[44512] = 32'hFFFFFFF1;
    // rom_array[44513] = 32'hFFFFFFF1;
    // rom_array[44514] = 32'hFFFFFFF1;
    // rom_array[44515] = 32'hFFFFFFF1;
    // rom_array[44516] = 32'hFFFFFFF1;
    // rom_array[44517] = 32'hFFFFFFF1;
    // rom_array[44518] = 32'hFFFFFFF1;
    // rom_array[44519] = 32'hFFFFFFF1;
    // rom_array[44520] = 32'hFFFFFFF1;
    // rom_array[44521] = 32'hFFFFFFF1;
    // rom_array[44522] = 32'hFFFFFFF1;
    // rom_array[44523] = 32'hFFFFFFF1;
    // rom_array[44524] = 32'hFFFFFFF1;
    // rom_array[44525] = 32'hFFFFFFF0;
    // rom_array[44526] = 32'hFFFFFFF0;
    // rom_array[44527] = 32'hFFFFFFF0;
    // rom_array[44528] = 32'hFFFFFFF0;
    // rom_array[44529] = 32'hFFFFFFF1;
    // rom_array[44530] = 32'hFFFFFFF1;
    // rom_array[44531] = 32'hFFFFFFF1;
    // rom_array[44532] = 32'hFFFFFFF1;
    // rom_array[44533] = 32'hFFFFFFF0;
    // rom_array[44534] = 32'hFFFFFFF0;
    // rom_array[44535] = 32'hFFFFFFF0;
    // rom_array[44536] = 32'hFFFFFFF0;
    // rom_array[44537] = 32'hFFFFFFF1;
    // rom_array[44538] = 32'hFFFFFFF1;
    // rom_array[44539] = 32'hFFFFFFF1;
    // rom_array[44540] = 32'hFFFFFFF1;
    // rom_array[44541] = 32'hFFFFFFF0;
    // rom_array[44542] = 32'hFFFFFFF0;
    // rom_array[44543] = 32'hFFFFFFF0;
    // rom_array[44544] = 32'hFFFFFFF0;
    // rom_array[44545] = 32'hFFFFFFF1;
    // rom_array[44546] = 32'hFFFFFFF1;
    // rom_array[44547] = 32'hFFFFFFF1;
    // rom_array[44548] = 32'hFFFFFFF1;
    // rom_array[44549] = 32'hFFFFFFF0;
    // rom_array[44550] = 32'hFFFFFFF0;
    // rom_array[44551] = 32'hFFFFFFF0;
    // rom_array[44552] = 32'hFFFFFFF0;
    // rom_array[44553] = 32'hFFFFFFF1;
    // rom_array[44554] = 32'hFFFFFFF1;
    // rom_array[44555] = 32'hFFFFFFF1;
    // rom_array[44556] = 32'hFFFFFFF1;
    // rom_array[44557] = 32'hFFFFFFF1;
    // rom_array[44558] = 32'hFFFFFFF1;
    // rom_array[44559] = 32'hFFFFFFF1;
    // rom_array[44560] = 32'hFFFFFFF1;
    // rom_array[44561] = 32'hFFFFFFF1;
    // rom_array[44562] = 32'hFFFFFFF1;
    // rom_array[44563] = 32'hFFFFFFF1;
    // rom_array[44564] = 32'hFFFFFFF1;
    // rom_array[44565] = 32'hFFFFFFF1;
    // rom_array[44566] = 32'hFFFFFFF1;
    // rom_array[44567] = 32'hFFFFFFF1;
    // rom_array[44568] = 32'hFFFFFFF1;
    // rom_array[44569] = 32'hFFFFFFF1;
    // rom_array[44570] = 32'hFFFFFFF1;
    // rom_array[44571] = 32'hFFFFFFF1;
    // rom_array[44572] = 32'hFFFFFFF1;
    // rom_array[44573] = 32'hFFFFFFF0;
    // rom_array[44574] = 32'hFFFFFFF0;
    // rom_array[44575] = 32'hFFFFFFF0;
    // rom_array[44576] = 32'hFFFFFFF0;
    // rom_array[44577] = 32'hFFFFFFF1;
    // rom_array[44578] = 32'hFFFFFFF1;
    // rom_array[44579] = 32'hFFFFFFF1;
    // rom_array[44580] = 32'hFFFFFFF1;
    // rom_array[44581] = 32'hFFFFFFF0;
    // rom_array[44582] = 32'hFFFFFFF0;
    // rom_array[44583] = 32'hFFFFFFF0;
    // rom_array[44584] = 32'hFFFFFFF0;
    // rom_array[44585] = 32'hFFFFFFF0;
    // rom_array[44586] = 32'hFFFFFFF0;
    // rom_array[44587] = 32'hFFFFFFF0;
    // rom_array[44588] = 32'hFFFFFFF0;
    // rom_array[44589] = 32'hFFFFFFF1;
    // rom_array[44590] = 32'hFFFFFFF1;
    // rom_array[44591] = 32'hFFFFFFF1;
    // rom_array[44592] = 32'hFFFFFFF1;
    // rom_array[44593] = 32'hFFFFFFF0;
    // rom_array[44594] = 32'hFFFFFFF0;
    // rom_array[44595] = 32'hFFFFFFF0;
    // rom_array[44596] = 32'hFFFFFFF0;
    // rom_array[44597] = 32'hFFFFFFF1;
    // rom_array[44598] = 32'hFFFFFFF1;
    // rom_array[44599] = 32'hFFFFFFF1;
    // rom_array[44600] = 32'hFFFFFFF1;
    // rom_array[44601] = 32'hFFFFFFF0;
    // rom_array[44602] = 32'hFFFFFFF0;
    // rom_array[44603] = 32'hFFFFFFF0;
    // rom_array[44604] = 32'hFFFFFFF0;
    // rom_array[44605] = 32'hFFFFFFF1;
    // rom_array[44606] = 32'hFFFFFFF1;
    // rom_array[44607] = 32'hFFFFFFF1;
    // rom_array[44608] = 32'hFFFFFFF1;
    // rom_array[44609] = 32'hFFFFFFF0;
    // rom_array[44610] = 32'hFFFFFFF0;
    // rom_array[44611] = 32'hFFFFFFF0;
    // rom_array[44612] = 32'hFFFFFFF0;
    // rom_array[44613] = 32'hFFFFFFF1;
    // rom_array[44614] = 32'hFFFFFFF1;
    // rom_array[44615] = 32'hFFFFFFF1;
    // rom_array[44616] = 32'hFFFFFFF1;
    // rom_array[44617] = 32'hFFFFFFF0;
    // rom_array[44618] = 32'hFFFFFFF0;
    // rom_array[44619] = 32'hFFFFFFF0;
    // rom_array[44620] = 32'hFFFFFFF0;
    // rom_array[44621] = 32'hFFFFFFF1;
    // rom_array[44622] = 32'hFFFFFFF1;
    // rom_array[44623] = 32'hFFFFFFF1;
    // rom_array[44624] = 32'hFFFFFFF1;
    // rom_array[44625] = 32'hFFFFFFF0;
    // rom_array[44626] = 32'hFFFFFFF0;
    // rom_array[44627] = 32'hFFFFFFF0;
    // rom_array[44628] = 32'hFFFFFFF0;
    // rom_array[44629] = 32'hFFFFFFF1;
    // rom_array[44630] = 32'hFFFFFFF1;
    // rom_array[44631] = 32'hFFFFFFF1;
    // rom_array[44632] = 32'hFFFFFFF1;
    // rom_array[44633] = 32'hFFFFFFF0;
    // rom_array[44634] = 32'hFFFFFFF0;
    // rom_array[44635] = 32'hFFFFFFF0;
    // rom_array[44636] = 32'hFFFFFFF0;
    // rom_array[44637] = 32'hFFFFFFF1;
    // rom_array[44638] = 32'hFFFFFFF1;
    // rom_array[44639] = 32'hFFFFFFF1;
    // rom_array[44640] = 32'hFFFFFFF1;
    // rom_array[44641] = 32'hFFFFFFF0;
    // rom_array[44642] = 32'hFFFFFFF0;
    // rom_array[44643] = 32'hFFFFFFF0;
    // rom_array[44644] = 32'hFFFFFFF0;
    // rom_array[44645] = 32'hFFFFFFF1;
    // rom_array[44646] = 32'hFFFFFFF1;
    // rom_array[44647] = 32'hFFFFFFF1;
    // rom_array[44648] = 32'hFFFFFFF1;
    // rom_array[44649] = 32'hFFFFFFF0;
    // rom_array[44650] = 32'hFFFFFFF0;
    // rom_array[44651] = 32'hFFFFFFF0;
    // rom_array[44652] = 32'hFFFFFFF0;
    // rom_array[44653] = 32'hFFFFFFF1;
    // rom_array[44654] = 32'hFFFFFFF1;
    // rom_array[44655] = 32'hFFFFFFF1;
    // rom_array[44656] = 32'hFFFFFFF1;
    // rom_array[44657] = 32'hFFFFFFF0;
    // rom_array[44658] = 32'hFFFFFFF0;
    // rom_array[44659] = 32'hFFFFFFF0;
    // rom_array[44660] = 32'hFFFFFFF0;
    // rom_array[44661] = 32'hFFFFFFF1;
    // rom_array[44662] = 32'hFFFFFFF1;
    // rom_array[44663] = 32'hFFFFFFF1;
    // rom_array[44664] = 32'hFFFFFFF1;
    // rom_array[44665] = 32'hFFFFFFF0;
    // rom_array[44666] = 32'hFFFFFFF0;
    // rom_array[44667] = 32'hFFFFFFF0;
    // rom_array[44668] = 32'hFFFFFFF0;
    // rom_array[44669] = 32'hFFFFFFF1;
    // rom_array[44670] = 32'hFFFFFFF1;
    // rom_array[44671] = 32'hFFFFFFF1;
    // rom_array[44672] = 32'hFFFFFFF1;
    // rom_array[44673] = 32'hFFFFFFF0;
    // rom_array[44674] = 32'hFFFFFFF0;
    // rom_array[44675] = 32'hFFFFFFF0;
    // rom_array[44676] = 32'hFFFFFFF0;
    // rom_array[44677] = 32'hFFFFFFF1;
    // rom_array[44678] = 32'hFFFFFFF1;
    // rom_array[44679] = 32'hFFFFFFF1;
    // rom_array[44680] = 32'hFFFFFFF1;
    // rom_array[44681] = 32'hFFFFFFF0;
    // rom_array[44682] = 32'hFFFFFFF0;
    // rom_array[44683] = 32'hFFFFFFF0;
    // rom_array[44684] = 32'hFFFFFFF0;
    // rom_array[44685] = 32'hFFFFFFF1;
    // rom_array[44686] = 32'hFFFFFFF1;
    // rom_array[44687] = 32'hFFFFFFF1;
    // rom_array[44688] = 32'hFFFFFFF1;
    // rom_array[44689] = 32'hFFFFFFF0;
    // rom_array[44690] = 32'hFFFFFFF0;
    // rom_array[44691] = 32'hFFFFFFF0;
    // rom_array[44692] = 32'hFFFFFFF0;
    // rom_array[44693] = 32'hFFFFFFF1;
    // rom_array[44694] = 32'hFFFFFFF1;
    // rom_array[44695] = 32'hFFFFFFF1;
    // rom_array[44696] = 32'hFFFFFFF1;
    // rom_array[44697] = 32'hFFFFFFF0;
    // rom_array[44698] = 32'hFFFFFFF0;
    // rom_array[44699] = 32'hFFFFFFF0;
    // rom_array[44700] = 32'hFFFFFFF0;
    // rom_array[44701] = 32'hFFFFFFF1;
    // rom_array[44702] = 32'hFFFFFFF1;
    // rom_array[44703] = 32'hFFFFFFF1;
    // rom_array[44704] = 32'hFFFFFFF1;
    // rom_array[44705] = 32'hFFFFFFF0;
    // rom_array[44706] = 32'hFFFFFFF0;
    // rom_array[44707] = 32'hFFFFFFF0;
    // rom_array[44708] = 32'hFFFFFFF0;
    // rom_array[44709] = 32'hFFFFFFF1;
    // rom_array[44710] = 32'hFFFFFFF1;
    // rom_array[44711] = 32'hFFFFFFF1;
    // rom_array[44712] = 32'hFFFFFFF1;
    // rom_array[44713] = 32'hFFFFFFF0;
    // rom_array[44714] = 32'hFFFFFFF0;
    // rom_array[44715] = 32'hFFFFFFF0;
    // rom_array[44716] = 32'hFFFFFFF0;
    // rom_array[44717] = 32'hFFFFFFF1;
    // rom_array[44718] = 32'hFFFFFFF1;
    // rom_array[44719] = 32'hFFFFFFF1;
    // rom_array[44720] = 32'hFFFFFFF1;
    // rom_array[44721] = 32'hFFFFFFF0;
    // rom_array[44722] = 32'hFFFFFFF0;
    // rom_array[44723] = 32'hFFFFFFF0;
    // rom_array[44724] = 32'hFFFFFFF0;
    // rom_array[44725] = 32'hFFFFFFF1;
    // rom_array[44726] = 32'hFFFFFFF1;
    // rom_array[44727] = 32'hFFFFFFF1;
    // rom_array[44728] = 32'hFFFFFFF1;
    // rom_array[44729] = 32'hFFFFFFF0;
    // rom_array[44730] = 32'hFFFFFFF0;
    // rom_array[44731] = 32'hFFFFFFF0;
    // rom_array[44732] = 32'hFFFFFFF0;
    // rom_array[44733] = 32'hFFFFFFF1;
    // rom_array[44734] = 32'hFFFFFFF1;
    // rom_array[44735] = 32'hFFFFFFF1;
    // rom_array[44736] = 32'hFFFFFFF1;
    // rom_array[44737] = 32'hFFFFFFF0;
    // rom_array[44738] = 32'hFFFFFFF0;
    // rom_array[44739] = 32'hFFFFFFF0;
    // rom_array[44740] = 32'hFFFFFFF0;
    // rom_array[44741] = 32'hFFFFFFF1;
    // rom_array[44742] = 32'hFFFFFFF1;
    // rom_array[44743] = 32'hFFFFFFF1;
    // rom_array[44744] = 32'hFFFFFFF1;
    // rom_array[44745] = 32'hFFFFFFF0;
    // rom_array[44746] = 32'hFFFFFFF0;
    // rom_array[44747] = 32'hFFFFFFF0;
    // rom_array[44748] = 32'hFFFFFFF0;
    // rom_array[44749] = 32'hFFFFFFF1;
    // rom_array[44750] = 32'hFFFFFFF1;
    // rom_array[44751] = 32'hFFFFFFF1;
    // rom_array[44752] = 32'hFFFFFFF1;
    // rom_array[44753] = 32'hFFFFFFF0;
    // rom_array[44754] = 32'hFFFFFFF0;
    // rom_array[44755] = 32'hFFFFFFF0;
    // rom_array[44756] = 32'hFFFFFFF0;
    // rom_array[44757] = 32'hFFFFFFF1;
    // rom_array[44758] = 32'hFFFFFFF1;
    // rom_array[44759] = 32'hFFFFFFF1;
    // rom_array[44760] = 32'hFFFFFFF1;
    // rom_array[44761] = 32'hFFFFFFF1;
    // rom_array[44762] = 32'hFFFFFFF1;
    // rom_array[44763] = 32'hFFFFFFF1;
    // rom_array[44764] = 32'hFFFFFFF1;
    // rom_array[44765] = 32'hFFFFFFF1;
    // rom_array[44766] = 32'hFFFFFFF1;
    // rom_array[44767] = 32'hFFFFFFF1;
    // rom_array[44768] = 32'hFFFFFFF1;
    // rom_array[44769] = 32'hFFFFFFF1;
    // rom_array[44770] = 32'hFFFFFFF1;
    // rom_array[44771] = 32'hFFFFFFF1;
    // rom_array[44772] = 32'hFFFFFFF1;
    // rom_array[44773] = 32'hFFFFFFF1;
    // rom_array[44774] = 32'hFFFFFFF1;
    // rom_array[44775] = 32'hFFFFFFF1;
    // rom_array[44776] = 32'hFFFFFFF1;
    // rom_array[44777] = 32'hFFFFFFF1;
    // rom_array[44778] = 32'hFFFFFFF1;
    // rom_array[44779] = 32'hFFFFFFF1;
    // rom_array[44780] = 32'hFFFFFFF1;
    // rom_array[44781] = 32'hFFFFFFF1;
    // rom_array[44782] = 32'hFFFFFFF1;
    // rom_array[44783] = 32'hFFFFFFF1;
    // rom_array[44784] = 32'hFFFFFFF1;
    // rom_array[44785] = 32'hFFFFFFF1;
    // rom_array[44786] = 32'hFFFFFFF1;
    // rom_array[44787] = 32'hFFFFFFF1;
    // rom_array[44788] = 32'hFFFFFFF1;
    // rom_array[44789] = 32'hFFFFFFF1;
    // rom_array[44790] = 32'hFFFFFFF1;
    // rom_array[44791] = 32'hFFFFFFF1;
    // rom_array[44792] = 32'hFFFFFFF1;
    // rom_array[44793] = 32'hFFFFFFF1;
    // rom_array[44794] = 32'hFFFFFFF1;
    // rom_array[44795] = 32'hFFFFFFF1;
    // rom_array[44796] = 32'hFFFFFFF1;
    // rom_array[44797] = 32'hFFFFFFF1;
    // rom_array[44798] = 32'hFFFFFFF1;
    // rom_array[44799] = 32'hFFFFFFF1;
    // rom_array[44800] = 32'hFFFFFFF1;
    // rom_array[44801] = 32'hFFFFFFF1;
    // rom_array[44802] = 32'hFFFFFFF1;
    // rom_array[44803] = 32'hFFFFFFF1;
    // rom_array[44804] = 32'hFFFFFFF1;
    // rom_array[44805] = 32'hFFFFFFF1;
    // rom_array[44806] = 32'hFFFFFFF1;
    // rom_array[44807] = 32'hFFFFFFF1;
    // rom_array[44808] = 32'hFFFFFFF1;
    // rom_array[44809] = 32'hFFFFFFF1;
    // rom_array[44810] = 32'hFFFFFFF1;
    // rom_array[44811] = 32'hFFFFFFF1;
    // rom_array[44812] = 32'hFFFFFFF1;
    // rom_array[44813] = 32'hFFFFFFF1;
    // rom_array[44814] = 32'hFFFFFFF1;
    // rom_array[44815] = 32'hFFFFFFF1;
    // rom_array[44816] = 32'hFFFFFFF1;
    // rom_array[44817] = 32'hFFFFFFF1;
    // rom_array[44818] = 32'hFFFFFFF1;
    // rom_array[44819] = 32'hFFFFFFF1;
    // rom_array[44820] = 32'hFFFFFFF1;
    // rom_array[44821] = 32'hFFFFFFF1;
    // rom_array[44822] = 32'hFFFFFFF1;
    // rom_array[44823] = 32'hFFFFFFF1;
    // rom_array[44824] = 32'hFFFFFFF1;
    // rom_array[44825] = 32'hFFFFFFF1;
    // rom_array[44826] = 32'hFFFFFFF1;
    // rom_array[44827] = 32'hFFFFFFF1;
    // rom_array[44828] = 32'hFFFFFFF1;
    // rom_array[44829] = 32'hFFFFFFF1;
    // rom_array[44830] = 32'hFFFFFFF1;
    // rom_array[44831] = 32'hFFFFFFF1;
    // rom_array[44832] = 32'hFFFFFFF1;
    // rom_array[44833] = 32'hFFFFFFF1;
    // rom_array[44834] = 32'hFFFFFFF1;
    // rom_array[44835] = 32'hFFFFFFF1;
    // rom_array[44836] = 32'hFFFFFFF1;
    // rom_array[44837] = 32'hFFFFFFF1;
    // rom_array[44838] = 32'hFFFFFFF1;
    // rom_array[44839] = 32'hFFFFFFF1;
    // rom_array[44840] = 32'hFFFFFFF1;
    // rom_array[44841] = 32'hFFFFFFF1;
    // rom_array[44842] = 32'hFFFFFFF1;
    // rom_array[44843] = 32'hFFFFFFF1;
    // rom_array[44844] = 32'hFFFFFFF1;
    // rom_array[44845] = 32'hFFFFFFF1;
    // rom_array[44846] = 32'hFFFFFFF1;
    // rom_array[44847] = 32'hFFFFFFF1;
    // rom_array[44848] = 32'hFFFFFFF1;
    // rom_array[44849] = 32'hFFFFFFF1;
    // rom_array[44850] = 32'hFFFFFFF1;
    // rom_array[44851] = 32'hFFFFFFF1;
    // rom_array[44852] = 32'hFFFFFFF1;
    // rom_array[44853] = 32'hFFFFFFF1;
    // rom_array[44854] = 32'hFFFFFFF1;
    // rom_array[44855] = 32'hFFFFFFF1;
    // rom_array[44856] = 32'hFFFFFFF1;
    // rom_array[44857] = 32'hFFFFFFF1;
    // rom_array[44858] = 32'hFFFFFFF1;
    // rom_array[44859] = 32'hFFFFFFF1;
    // rom_array[44860] = 32'hFFFFFFF1;
    // rom_array[44861] = 32'hFFFFFFF1;
    // rom_array[44862] = 32'hFFFFFFF1;
    // rom_array[44863] = 32'hFFFFFFF1;
    // rom_array[44864] = 32'hFFFFFFF1;
    // rom_array[44865] = 32'hFFFFFFF1;
    // rom_array[44866] = 32'hFFFFFFF1;
    // rom_array[44867] = 32'hFFFFFFF1;
    // rom_array[44868] = 32'hFFFFFFF1;
    // rom_array[44869] = 32'hFFFFFFF1;
    // rom_array[44870] = 32'hFFFFFFF1;
    // rom_array[44871] = 32'hFFFFFFF1;
    // rom_array[44872] = 32'hFFFFFFF1;
    // rom_array[44873] = 32'hFFFFFFF0;
    // rom_array[44874] = 32'hFFFFFFF0;
    // rom_array[44875] = 32'hFFFFFFF0;
    // rom_array[44876] = 32'hFFFFFFF0;
    // rom_array[44877] = 32'hFFFFFFF1;
    // rom_array[44878] = 32'hFFFFFFF1;
    // rom_array[44879] = 32'hFFFFFFF1;
    // rom_array[44880] = 32'hFFFFFFF1;
    // rom_array[44881] = 32'hFFFFFFF0;
    // rom_array[44882] = 32'hFFFFFFF0;
    // rom_array[44883] = 32'hFFFFFFF0;
    // rom_array[44884] = 32'hFFFFFFF0;
    // rom_array[44885] = 32'hFFFFFFF1;
    // rom_array[44886] = 32'hFFFFFFF1;
    // rom_array[44887] = 32'hFFFFFFF1;
    // rom_array[44888] = 32'hFFFFFFF1;
    // rom_array[44889] = 32'hFFFFFFF0;
    // rom_array[44890] = 32'hFFFFFFF0;
    // rom_array[44891] = 32'hFFFFFFF0;
    // rom_array[44892] = 32'hFFFFFFF0;
    // rom_array[44893] = 32'hFFFFFFF1;
    // rom_array[44894] = 32'hFFFFFFF1;
    // rom_array[44895] = 32'hFFFFFFF1;
    // rom_array[44896] = 32'hFFFFFFF1;
    // rom_array[44897] = 32'hFFFFFFF0;
    // rom_array[44898] = 32'hFFFFFFF0;
    // rom_array[44899] = 32'hFFFFFFF0;
    // rom_array[44900] = 32'hFFFFFFF0;
    // rom_array[44901] = 32'hFFFFFFF1;
    // rom_array[44902] = 32'hFFFFFFF1;
    // rom_array[44903] = 32'hFFFFFFF1;
    // rom_array[44904] = 32'hFFFFFFF1;
    // rom_array[44905] = 32'hFFFFFFF0;
    // rom_array[44906] = 32'hFFFFFFF0;
    // rom_array[44907] = 32'hFFFFFFF0;
    // rom_array[44908] = 32'hFFFFFFF0;
    // rom_array[44909] = 32'hFFFFFFF1;
    // rom_array[44910] = 32'hFFFFFFF1;
    // rom_array[44911] = 32'hFFFFFFF1;
    // rom_array[44912] = 32'hFFFFFFF1;
    // rom_array[44913] = 32'hFFFFFFF0;
    // rom_array[44914] = 32'hFFFFFFF0;
    // rom_array[44915] = 32'hFFFFFFF0;
    // rom_array[44916] = 32'hFFFFFFF0;
    // rom_array[44917] = 32'hFFFFFFF1;
    // rom_array[44918] = 32'hFFFFFFF1;
    // rom_array[44919] = 32'hFFFFFFF1;
    // rom_array[44920] = 32'hFFFFFFF1;
    // rom_array[44921] = 32'hFFFFFFF0;
    // rom_array[44922] = 32'hFFFFFFF0;
    // rom_array[44923] = 32'hFFFFFFF0;
    // rom_array[44924] = 32'hFFFFFFF0;
    // rom_array[44925] = 32'hFFFFFFF1;
    // rom_array[44926] = 32'hFFFFFFF1;
    // rom_array[44927] = 32'hFFFFFFF1;
    // rom_array[44928] = 32'hFFFFFFF1;
    // rom_array[44929] = 32'hFFFFFFF0;
    // rom_array[44930] = 32'hFFFFFFF0;
    // rom_array[44931] = 32'hFFFFFFF0;
    // rom_array[44932] = 32'hFFFFFFF0;
    // rom_array[44933] = 32'hFFFFFFF1;
    // rom_array[44934] = 32'hFFFFFFF1;
    // rom_array[44935] = 32'hFFFFFFF1;
    // rom_array[44936] = 32'hFFFFFFF1;
    // rom_array[44937] = 32'hFFFFFFF0;
    // rom_array[44938] = 32'hFFFFFFF0;
    // rom_array[44939] = 32'hFFFFFFF0;
    // rom_array[44940] = 32'hFFFFFFF0;
    // rom_array[44941] = 32'hFFFFFFF1;
    // rom_array[44942] = 32'hFFFFFFF1;
    // rom_array[44943] = 32'hFFFFFFF1;
    // rom_array[44944] = 32'hFFFFFFF1;
    // rom_array[44945] = 32'hFFFFFFF0;
    // rom_array[44946] = 32'hFFFFFFF0;
    // rom_array[44947] = 32'hFFFFFFF0;
    // rom_array[44948] = 32'hFFFFFFF0;
    // rom_array[44949] = 32'hFFFFFFF1;
    // rom_array[44950] = 32'hFFFFFFF1;
    // rom_array[44951] = 32'hFFFFFFF1;
    // rom_array[44952] = 32'hFFFFFFF1;
    // rom_array[44953] = 32'hFFFFFFF0;
    // rom_array[44954] = 32'hFFFFFFF0;
    // rom_array[44955] = 32'hFFFFFFF0;
    // rom_array[44956] = 32'hFFFFFFF0;
    // rom_array[44957] = 32'hFFFFFFF1;
    // rom_array[44958] = 32'hFFFFFFF1;
    // rom_array[44959] = 32'hFFFFFFF1;
    // rom_array[44960] = 32'hFFFFFFF1;
    // rom_array[44961] = 32'hFFFFFFF0;
    // rom_array[44962] = 32'hFFFFFFF0;
    // rom_array[44963] = 32'hFFFFFFF0;
    // rom_array[44964] = 32'hFFFFFFF0;
    // rom_array[44965] = 32'hFFFFFFF1;
    // rom_array[44966] = 32'hFFFFFFF1;
    // rom_array[44967] = 32'hFFFFFFF1;
    // rom_array[44968] = 32'hFFFFFFF1;
    // rom_array[44969] = 32'hFFFFFFF0;
    // rom_array[44970] = 32'hFFFFFFF0;
    // rom_array[44971] = 32'hFFFFFFF0;
    // rom_array[44972] = 32'hFFFFFFF0;
    // rom_array[44973] = 32'hFFFFFFF1;
    // rom_array[44974] = 32'hFFFFFFF1;
    // rom_array[44975] = 32'hFFFFFFF1;
    // rom_array[44976] = 32'hFFFFFFF1;
    // rom_array[44977] = 32'hFFFFFFF0;
    // rom_array[44978] = 32'hFFFFFFF0;
    // rom_array[44979] = 32'hFFFFFFF0;
    // rom_array[44980] = 32'hFFFFFFF0;
    // rom_array[44981] = 32'hFFFFFFF1;
    // rom_array[44982] = 32'hFFFFFFF1;
    // rom_array[44983] = 32'hFFFFFFF1;
    // rom_array[44984] = 32'hFFFFFFF1;
    // rom_array[44985] = 32'hFFFFFFF0;
    // rom_array[44986] = 32'hFFFFFFF0;
    // rom_array[44987] = 32'hFFFFFFF0;
    // rom_array[44988] = 32'hFFFFFFF0;
    // rom_array[44989] = 32'hFFFFFFF1;
    // rom_array[44990] = 32'hFFFFFFF1;
    // rom_array[44991] = 32'hFFFFFFF1;
    // rom_array[44992] = 32'hFFFFFFF1;
    // rom_array[44993] = 32'hFFFFFFF0;
    // rom_array[44994] = 32'hFFFFFFF0;
    // rom_array[44995] = 32'hFFFFFFF0;
    // rom_array[44996] = 32'hFFFFFFF0;
    // rom_array[44997] = 32'hFFFFFFF1;
    // rom_array[44998] = 32'hFFFFFFF1;
    // rom_array[44999] = 32'hFFFFFFF1;
    // rom_array[45000] = 32'hFFFFFFF1;
    // rom_array[45001] = 32'hFFFFFFF0;
    // rom_array[45002] = 32'hFFFFFFF0;
    // rom_array[45003] = 32'hFFFFFFF1;
    // rom_array[45004] = 32'hFFFFFFF1;
    // rom_array[45005] = 32'hFFFFFFF0;
    // rom_array[45006] = 32'hFFFFFFF0;
    // rom_array[45007] = 32'hFFFFFFF1;
    // rom_array[45008] = 32'hFFFFFFF1;
    // rom_array[45009] = 32'hFFFFFFF0;
    // rom_array[45010] = 32'hFFFFFFF0;
    // rom_array[45011] = 32'hFFFFFFF1;
    // rom_array[45012] = 32'hFFFFFFF1;
    // rom_array[45013] = 32'hFFFFFFF0;
    // rom_array[45014] = 32'hFFFFFFF0;
    // rom_array[45015] = 32'hFFFFFFF1;
    // rom_array[45016] = 32'hFFFFFFF1;
    // rom_array[45017] = 32'hFFFFFFF0;
    // rom_array[45018] = 32'hFFFFFFF0;
    // rom_array[45019] = 32'hFFFFFFF1;
    // rom_array[45020] = 32'hFFFFFFF1;
    // rom_array[45021] = 32'hFFFFFFF0;
    // rom_array[45022] = 32'hFFFFFFF0;
    // rom_array[45023] = 32'hFFFFFFF1;
    // rom_array[45024] = 32'hFFFFFFF1;
    // rom_array[45025] = 32'hFFFFFFF0;
    // rom_array[45026] = 32'hFFFFFFF0;
    // rom_array[45027] = 32'hFFFFFFF1;
    // rom_array[45028] = 32'hFFFFFFF1;
    // rom_array[45029] = 32'hFFFFFFF0;
    // rom_array[45030] = 32'hFFFFFFF0;
    // rom_array[45031] = 32'hFFFFFFF1;
    // rom_array[45032] = 32'hFFFFFFF1;
    // rom_array[45033] = 32'hFFFFFFF0;
    // rom_array[45034] = 32'hFFFFFFF0;
    // rom_array[45035] = 32'hFFFFFFF1;
    // rom_array[45036] = 32'hFFFFFFF1;
    // rom_array[45037] = 32'hFFFFFFF0;
    // rom_array[45038] = 32'hFFFFFFF0;
    // rom_array[45039] = 32'hFFFFFFF1;
    // rom_array[45040] = 32'hFFFFFFF1;
    // rom_array[45041] = 32'hFFFFFFF0;
    // rom_array[45042] = 32'hFFFFFFF0;
    // rom_array[45043] = 32'hFFFFFFF1;
    // rom_array[45044] = 32'hFFFFFFF1;
    // rom_array[45045] = 32'hFFFFFFF0;
    // rom_array[45046] = 32'hFFFFFFF0;
    // rom_array[45047] = 32'hFFFFFFF1;
    // rom_array[45048] = 32'hFFFFFFF1;
    // rom_array[45049] = 32'hFFFFFFF1;
    // rom_array[45050] = 32'hFFFFFFF1;
    // rom_array[45051] = 32'hFFFFFFF1;
    // rom_array[45052] = 32'hFFFFFFF1;
    // rom_array[45053] = 32'hFFFFFFF0;
    // rom_array[45054] = 32'hFFFFFFF0;
    // rom_array[45055] = 32'hFFFFFFF0;
    // rom_array[45056] = 32'hFFFFFFF0;
    // rom_array[45057] = 32'hFFFFFFF1;
    // rom_array[45058] = 32'hFFFFFFF1;
    // rom_array[45059] = 32'hFFFFFFF1;
    // rom_array[45060] = 32'hFFFFFFF1;
    // rom_array[45061] = 32'hFFFFFFF0;
    // rom_array[45062] = 32'hFFFFFFF0;
    // rom_array[45063] = 32'hFFFFFFF0;
    // rom_array[45064] = 32'hFFFFFFF0;
    // rom_array[45065] = 32'hFFFFFFF1;
    // rom_array[45066] = 32'hFFFFFFF1;
    // rom_array[45067] = 32'hFFFFFFF1;
    // rom_array[45068] = 32'hFFFFFFF1;
    // rom_array[45069] = 32'hFFFFFFF0;
    // rom_array[45070] = 32'hFFFFFFF0;
    // rom_array[45071] = 32'hFFFFFFF0;
    // rom_array[45072] = 32'hFFFFFFF0;
    // rom_array[45073] = 32'hFFFFFFF1;
    // rom_array[45074] = 32'hFFFFFFF1;
    // rom_array[45075] = 32'hFFFFFFF1;
    // rom_array[45076] = 32'hFFFFFFF1;
    // rom_array[45077] = 32'hFFFFFFF0;
    // rom_array[45078] = 32'hFFFFFFF0;
    // rom_array[45079] = 32'hFFFFFFF0;
    // rom_array[45080] = 32'hFFFFFFF0;
    // rom_array[45081] = 32'hFFFFFFF1;
    // rom_array[45082] = 32'hFFFFFFF1;
    // rom_array[45083] = 32'hFFFFFFF1;
    // rom_array[45084] = 32'hFFFFFFF1;
    // rom_array[45085] = 32'hFFFFFFF0;
    // rom_array[45086] = 32'hFFFFFFF0;
    // rom_array[45087] = 32'hFFFFFFF0;
    // rom_array[45088] = 32'hFFFFFFF0;
    // rom_array[45089] = 32'hFFFFFFF1;
    // rom_array[45090] = 32'hFFFFFFF1;
    // rom_array[45091] = 32'hFFFFFFF1;
    // rom_array[45092] = 32'hFFFFFFF1;
    // rom_array[45093] = 32'hFFFFFFF0;
    // rom_array[45094] = 32'hFFFFFFF0;
    // rom_array[45095] = 32'hFFFFFFF0;
    // rom_array[45096] = 32'hFFFFFFF0;
    // rom_array[45097] = 32'hFFFFFFF1;
    // rom_array[45098] = 32'hFFFFFFF1;
    // rom_array[45099] = 32'hFFFFFFF1;
    // rom_array[45100] = 32'hFFFFFFF1;
    // rom_array[45101] = 32'hFFFFFFF0;
    // rom_array[45102] = 32'hFFFFFFF0;
    // rom_array[45103] = 32'hFFFFFFF0;
    // rom_array[45104] = 32'hFFFFFFF0;
    // rom_array[45105] = 32'hFFFFFFF1;
    // rom_array[45106] = 32'hFFFFFFF1;
    // rom_array[45107] = 32'hFFFFFFF1;
    // rom_array[45108] = 32'hFFFFFFF1;
    // rom_array[45109] = 32'hFFFFFFF0;
    // rom_array[45110] = 32'hFFFFFFF0;
    // rom_array[45111] = 32'hFFFFFFF0;
    // rom_array[45112] = 32'hFFFFFFF0;
    // rom_array[45113] = 32'hFFFFFFF1;
    // rom_array[45114] = 32'hFFFFFFF1;
    // rom_array[45115] = 32'hFFFFFFF1;
    // rom_array[45116] = 32'hFFFFFFF1;
    // rom_array[45117] = 32'hFFFFFFF0;
    // rom_array[45118] = 32'hFFFFFFF0;
    // rom_array[45119] = 32'hFFFFFFF0;
    // rom_array[45120] = 32'hFFFFFFF0;
    // rom_array[45121] = 32'hFFFFFFF1;
    // rom_array[45122] = 32'hFFFFFFF1;
    // rom_array[45123] = 32'hFFFFFFF1;
    // rom_array[45124] = 32'hFFFFFFF1;
    // rom_array[45125] = 32'hFFFFFFF0;
    // rom_array[45126] = 32'hFFFFFFF0;
    // rom_array[45127] = 32'hFFFFFFF0;
    // rom_array[45128] = 32'hFFFFFFF0;
    // rom_array[45129] = 32'hFFFFFFF1;
    // rom_array[45130] = 32'hFFFFFFF1;
    // rom_array[45131] = 32'hFFFFFFF1;
    // rom_array[45132] = 32'hFFFFFFF1;
    // rom_array[45133] = 32'hFFFFFFF0;
    // rom_array[45134] = 32'hFFFFFFF0;
    // rom_array[45135] = 32'hFFFFFFF0;
    // rom_array[45136] = 32'hFFFFFFF0;
    // rom_array[45137] = 32'hFFFFFFF1;
    // rom_array[45138] = 32'hFFFFFFF1;
    // rom_array[45139] = 32'hFFFFFFF1;
    // rom_array[45140] = 32'hFFFFFFF1;
    // rom_array[45141] = 32'hFFFFFFF0;
    // rom_array[45142] = 32'hFFFFFFF0;
    // rom_array[45143] = 32'hFFFFFFF0;
    // rom_array[45144] = 32'hFFFFFFF0;
    // rom_array[45145] = 32'hFFFFFFF1;
    // rom_array[45146] = 32'hFFFFFFF1;
    // rom_array[45147] = 32'hFFFFFFF1;
    // rom_array[45148] = 32'hFFFFFFF1;
    // rom_array[45149] = 32'hFFFFFFF0;
    // rom_array[45150] = 32'hFFFFFFF0;
    // rom_array[45151] = 32'hFFFFFFF0;
    // rom_array[45152] = 32'hFFFFFFF0;
    // rom_array[45153] = 32'hFFFFFFF1;
    // rom_array[45154] = 32'hFFFFFFF1;
    // rom_array[45155] = 32'hFFFFFFF1;
    // rom_array[45156] = 32'hFFFFFFF1;
    // rom_array[45157] = 32'hFFFFFFF0;
    // rom_array[45158] = 32'hFFFFFFF0;
    // rom_array[45159] = 32'hFFFFFFF0;
    // rom_array[45160] = 32'hFFFFFFF0;
    // rom_array[45161] = 32'hFFFFFFF1;
    // rom_array[45162] = 32'hFFFFFFF1;
    // rom_array[45163] = 32'hFFFFFFF1;
    // rom_array[45164] = 32'hFFFFFFF1;
    // rom_array[45165] = 32'hFFFFFFF0;
    // rom_array[45166] = 32'hFFFFFFF0;
    // rom_array[45167] = 32'hFFFFFFF0;
    // rom_array[45168] = 32'hFFFFFFF0;
    // rom_array[45169] = 32'hFFFFFFF1;
    // rom_array[45170] = 32'hFFFFFFF1;
    // rom_array[45171] = 32'hFFFFFFF1;
    // rom_array[45172] = 32'hFFFFFFF1;
    // rom_array[45173] = 32'hFFFFFFF0;
    // rom_array[45174] = 32'hFFFFFFF0;
    // rom_array[45175] = 32'hFFFFFFF0;
    // rom_array[45176] = 32'hFFFFFFF0;
    // rom_array[45177] = 32'hFFFFFFF0;
    // rom_array[45178] = 32'hFFFFFFF0;
    // rom_array[45179] = 32'hFFFFFFF0;
    // rom_array[45180] = 32'hFFFFFFF0;
    // rom_array[45181] = 32'hFFFFFFF1;
    // rom_array[45182] = 32'hFFFFFFF1;
    // rom_array[45183] = 32'hFFFFFFF1;
    // rom_array[45184] = 32'hFFFFFFF1;
    // rom_array[45185] = 32'hFFFFFFF0;
    // rom_array[45186] = 32'hFFFFFFF0;
    // rom_array[45187] = 32'hFFFFFFF0;
    // rom_array[45188] = 32'hFFFFFFF0;
    // rom_array[45189] = 32'hFFFFFFF1;
    // rom_array[45190] = 32'hFFFFFFF1;
    // rom_array[45191] = 32'hFFFFFFF1;
    // rom_array[45192] = 32'hFFFFFFF1;
    // rom_array[45193] = 32'hFFFFFFF0;
    // rom_array[45194] = 32'hFFFFFFF0;
    // rom_array[45195] = 32'hFFFFFFF0;
    // rom_array[45196] = 32'hFFFFFFF0;
    // rom_array[45197] = 32'hFFFFFFF1;
    // rom_array[45198] = 32'hFFFFFFF1;
    // rom_array[45199] = 32'hFFFFFFF1;
    // rom_array[45200] = 32'hFFFFFFF1;
    // rom_array[45201] = 32'hFFFFFFF0;
    // rom_array[45202] = 32'hFFFFFFF0;
    // rom_array[45203] = 32'hFFFFFFF0;
    // rom_array[45204] = 32'hFFFFFFF0;
    // rom_array[45205] = 32'hFFFFFFF1;
    // rom_array[45206] = 32'hFFFFFFF1;
    // rom_array[45207] = 32'hFFFFFFF1;
    // rom_array[45208] = 32'hFFFFFFF1;
    // rom_array[45209] = 32'hFFFFFFF1;
    // rom_array[45210] = 32'hFFFFFFF1;
    // rom_array[45211] = 32'hFFFFFFF1;
    // rom_array[45212] = 32'hFFFFFFF1;
    // rom_array[45213] = 32'hFFFFFFF1;
    // rom_array[45214] = 32'hFFFFFFF1;
    // rom_array[45215] = 32'hFFFFFFF1;
    // rom_array[45216] = 32'hFFFFFFF1;
    // rom_array[45217] = 32'hFFFFFFF1;
    // rom_array[45218] = 32'hFFFFFFF1;
    // rom_array[45219] = 32'hFFFFFFF1;
    // rom_array[45220] = 32'hFFFFFFF1;
    // rom_array[45221] = 32'hFFFFFFF1;
    // rom_array[45222] = 32'hFFFFFFF1;
    // rom_array[45223] = 32'hFFFFFFF1;
    // rom_array[45224] = 32'hFFFFFFF1;
    // rom_array[45225] = 32'hFFFFFFF1;
    // rom_array[45226] = 32'hFFFFFFF1;
    // rom_array[45227] = 32'hFFFFFFF1;
    // rom_array[45228] = 32'hFFFFFFF1;
    // rom_array[45229] = 32'hFFFFFFF1;
    // rom_array[45230] = 32'hFFFFFFF1;
    // rom_array[45231] = 32'hFFFFFFF1;
    // rom_array[45232] = 32'hFFFFFFF1;
    // rom_array[45233] = 32'hFFFFFFF1;
    // rom_array[45234] = 32'hFFFFFFF1;
    // rom_array[45235] = 32'hFFFFFFF1;
    // rom_array[45236] = 32'hFFFFFFF1;
    // rom_array[45237] = 32'hFFFFFFF1;
    // rom_array[45238] = 32'hFFFFFFF1;
    // rom_array[45239] = 32'hFFFFFFF1;
    // rom_array[45240] = 32'hFFFFFFF1;
    // rom_array[45241] = 32'hFFFFFFF1;
    // rom_array[45242] = 32'hFFFFFFF1;
    // rom_array[45243] = 32'hFFFFFFF1;
    // rom_array[45244] = 32'hFFFFFFF1;
    // rom_array[45245] = 32'hFFFFFFF1;
    // rom_array[45246] = 32'hFFFFFFF1;
    // rom_array[45247] = 32'hFFFFFFF1;
    // rom_array[45248] = 32'hFFFFFFF1;
    // rom_array[45249] = 32'hFFFFFFF1;
    // rom_array[45250] = 32'hFFFFFFF1;
    // rom_array[45251] = 32'hFFFFFFF1;
    // rom_array[45252] = 32'hFFFFFFF1;
    // rom_array[45253] = 32'hFFFFFFF1;
    // rom_array[45254] = 32'hFFFFFFF1;
    // rom_array[45255] = 32'hFFFFFFF1;
    // rom_array[45256] = 32'hFFFFFFF1;
    // rom_array[45257] = 32'hFFFFFFF1;
    // rom_array[45258] = 32'hFFFFFFF1;
    // rom_array[45259] = 32'hFFFFFFF1;
    // rom_array[45260] = 32'hFFFFFFF1;
    // rom_array[45261] = 32'hFFFFFFF1;
    // rom_array[45262] = 32'hFFFFFFF1;
    // rom_array[45263] = 32'hFFFFFFF1;
    // rom_array[45264] = 32'hFFFFFFF1;
    // rom_array[45265] = 32'hFFFFFFF1;
    // rom_array[45266] = 32'hFFFFFFF1;
    // rom_array[45267] = 32'hFFFFFFF1;
    // rom_array[45268] = 32'hFFFFFFF1;
    // rom_array[45269] = 32'hFFFFFFF1;
    // rom_array[45270] = 32'hFFFFFFF1;
    // rom_array[45271] = 32'hFFFFFFF1;
    // rom_array[45272] = 32'hFFFFFFF1;
    // rom_array[45273] = 32'hFFFFFFF1;
    // rom_array[45274] = 32'hFFFFFFF1;
    // rom_array[45275] = 32'hFFFFFFF1;
    // rom_array[45276] = 32'hFFFFFFF1;
    // rom_array[45277] = 32'hFFFFFFF0;
    // rom_array[45278] = 32'hFFFFFFF0;
    // rom_array[45279] = 32'hFFFFFFF0;
    // rom_array[45280] = 32'hFFFFFFF0;
    // rom_array[45281] = 32'hFFFFFFF1;
    // rom_array[45282] = 32'hFFFFFFF1;
    // rom_array[45283] = 32'hFFFFFFF1;
    // rom_array[45284] = 32'hFFFFFFF1;
    // rom_array[45285] = 32'hFFFFFFF0;
    // rom_array[45286] = 32'hFFFFFFF0;
    // rom_array[45287] = 32'hFFFFFFF0;
    // rom_array[45288] = 32'hFFFFFFF0;
    // rom_array[45289] = 32'hFFFFFFF1;
    // rom_array[45290] = 32'hFFFFFFF1;
    // rom_array[45291] = 32'hFFFFFFF1;
    // rom_array[45292] = 32'hFFFFFFF1;
    // rom_array[45293] = 32'hFFFFFFF0;
    // rom_array[45294] = 32'hFFFFFFF0;
    // rom_array[45295] = 32'hFFFFFFF0;
    // rom_array[45296] = 32'hFFFFFFF0;
    // rom_array[45297] = 32'hFFFFFFF1;
    // rom_array[45298] = 32'hFFFFFFF1;
    // rom_array[45299] = 32'hFFFFFFF1;
    // rom_array[45300] = 32'hFFFFFFF1;
    // rom_array[45301] = 32'hFFFFFFF0;
    // rom_array[45302] = 32'hFFFFFFF0;
    // rom_array[45303] = 32'hFFFFFFF0;
    // rom_array[45304] = 32'hFFFFFFF0;
    // rom_array[45305] = 32'hFFFFFFF1;
    // rom_array[45306] = 32'hFFFFFFF1;
    // rom_array[45307] = 32'hFFFFFFF1;
    // rom_array[45308] = 32'hFFFFFFF1;
    // rom_array[45309] = 32'hFFFFFFF1;
    // rom_array[45310] = 32'hFFFFFFF1;
    // rom_array[45311] = 32'hFFFFFFF1;
    // rom_array[45312] = 32'hFFFFFFF1;
    // rom_array[45313] = 32'hFFFFFFF1;
    // rom_array[45314] = 32'hFFFFFFF1;
    // rom_array[45315] = 32'hFFFFFFF1;
    // rom_array[45316] = 32'hFFFFFFF1;
    // rom_array[45317] = 32'hFFFFFFF1;
    // rom_array[45318] = 32'hFFFFFFF1;
    // rom_array[45319] = 32'hFFFFFFF1;
    // rom_array[45320] = 32'hFFFFFFF1;
    // rom_array[45321] = 32'hFFFFFFF1;
    // rom_array[45322] = 32'hFFFFFFF1;
    // rom_array[45323] = 32'hFFFFFFF1;
    // rom_array[45324] = 32'hFFFFFFF1;
    // rom_array[45325] = 32'hFFFFFFF1;
    // rom_array[45326] = 32'hFFFFFFF1;
    // rom_array[45327] = 32'hFFFFFFF1;
    // rom_array[45328] = 32'hFFFFFFF1;
    // rom_array[45329] = 32'hFFFFFFF1;
    // rom_array[45330] = 32'hFFFFFFF1;
    // rom_array[45331] = 32'hFFFFFFF1;
    // rom_array[45332] = 32'hFFFFFFF1;
    // rom_array[45333] = 32'hFFFFFFF1;
    // rom_array[45334] = 32'hFFFFFFF1;
    // rom_array[45335] = 32'hFFFFFFF1;
    // rom_array[45336] = 32'hFFFFFFF1;
    // rom_array[45337] = 32'hFFFFFFF1;
    // rom_array[45338] = 32'hFFFFFFF1;
    // rom_array[45339] = 32'hFFFFFFF1;
    // rom_array[45340] = 32'hFFFFFFF1;
    // rom_array[45341] = 32'hFFFFFFF1;
    // rom_array[45342] = 32'hFFFFFFF1;
    // rom_array[45343] = 32'hFFFFFFF1;
    // rom_array[45344] = 32'hFFFFFFF1;
    // rom_array[45345] = 32'hFFFFFFF1;
    // rom_array[45346] = 32'hFFFFFFF1;
    // rom_array[45347] = 32'hFFFFFFF1;
    // rom_array[45348] = 32'hFFFFFFF1;
    // rom_array[45349] = 32'hFFFFFFF1;
    // rom_array[45350] = 32'hFFFFFFF1;
    // rom_array[45351] = 32'hFFFFFFF1;
    // rom_array[45352] = 32'hFFFFFFF1;
    // rom_array[45353] = 32'hFFFFFFF1;
    // rom_array[45354] = 32'hFFFFFFF1;
    // rom_array[45355] = 32'hFFFFFFF1;
    // rom_array[45356] = 32'hFFFFFFF1;
    // rom_array[45357] = 32'hFFFFFFF1;
    // rom_array[45358] = 32'hFFFFFFF1;
    // rom_array[45359] = 32'hFFFFFFF1;
    // rom_array[45360] = 32'hFFFFFFF1;
    // rom_array[45361] = 32'hFFFFFFF1;
    // rom_array[45362] = 32'hFFFFFFF1;
    // rom_array[45363] = 32'hFFFFFFF1;
    // rom_array[45364] = 32'hFFFFFFF1;
    // rom_array[45365] = 32'hFFFFFFF1;
    // rom_array[45366] = 32'hFFFFFFF1;
    // rom_array[45367] = 32'hFFFFFFF1;
    // rom_array[45368] = 32'hFFFFFFF1;
    // rom_array[45369] = 32'hFFFFFFF1;
    // rom_array[45370] = 32'hFFFFFFF1;
    // rom_array[45371] = 32'hFFFFFFF1;
    // rom_array[45372] = 32'hFFFFFFF1;
    // rom_array[45373] = 32'hFFFFFFF0;
    // rom_array[45374] = 32'hFFFFFFF0;
    // rom_array[45375] = 32'hFFFFFFF0;
    // rom_array[45376] = 32'hFFFFFFF0;
    // rom_array[45377] = 32'hFFFFFFF1;
    // rom_array[45378] = 32'hFFFFFFF1;
    // rom_array[45379] = 32'hFFFFFFF1;
    // rom_array[45380] = 32'hFFFFFFF1;
    // rom_array[45381] = 32'hFFFFFFF0;
    // rom_array[45382] = 32'hFFFFFFF0;
    // rom_array[45383] = 32'hFFFFFFF0;
    // rom_array[45384] = 32'hFFFFFFF0;
    // rom_array[45385] = 32'hFFFFFFF1;
    // rom_array[45386] = 32'hFFFFFFF1;
    // rom_array[45387] = 32'hFFFFFFF1;
    // rom_array[45388] = 32'hFFFFFFF1;
    // rom_array[45389] = 32'hFFFFFFF0;
    // rom_array[45390] = 32'hFFFFFFF0;
    // rom_array[45391] = 32'hFFFFFFF0;
    // rom_array[45392] = 32'hFFFFFFF0;
    // rom_array[45393] = 32'hFFFFFFF1;
    // rom_array[45394] = 32'hFFFFFFF1;
    // rom_array[45395] = 32'hFFFFFFF1;
    // rom_array[45396] = 32'hFFFFFFF1;
    // rom_array[45397] = 32'hFFFFFFF0;
    // rom_array[45398] = 32'hFFFFFFF0;
    // rom_array[45399] = 32'hFFFFFFF0;
    // rom_array[45400] = 32'hFFFFFFF0;
    // rom_array[45401] = 32'hFFFFFFF1;
    // rom_array[45402] = 32'hFFFFFFF1;
    // rom_array[45403] = 32'hFFFFFFF1;
    // rom_array[45404] = 32'hFFFFFFF1;
    // rom_array[45405] = 32'hFFFFFFF0;
    // rom_array[45406] = 32'hFFFFFFF0;
    // rom_array[45407] = 32'hFFFFFFF0;
    // rom_array[45408] = 32'hFFFFFFF0;
    // rom_array[45409] = 32'hFFFFFFF1;
    // rom_array[45410] = 32'hFFFFFFF1;
    // rom_array[45411] = 32'hFFFFFFF1;
    // rom_array[45412] = 32'hFFFFFFF1;
    // rom_array[45413] = 32'hFFFFFFF0;
    // rom_array[45414] = 32'hFFFFFFF0;
    // rom_array[45415] = 32'hFFFFFFF0;
    // rom_array[45416] = 32'hFFFFFFF0;
    // rom_array[45417] = 32'hFFFFFFF1;
    // rom_array[45418] = 32'hFFFFFFF1;
    // rom_array[45419] = 32'hFFFFFFF1;
    // rom_array[45420] = 32'hFFFFFFF1;
    // rom_array[45421] = 32'hFFFFFFF0;
    // rom_array[45422] = 32'hFFFFFFF0;
    // rom_array[45423] = 32'hFFFFFFF0;
    // rom_array[45424] = 32'hFFFFFFF0;
    // rom_array[45425] = 32'hFFFFFFF1;
    // rom_array[45426] = 32'hFFFFFFF1;
    // rom_array[45427] = 32'hFFFFFFF1;
    // rom_array[45428] = 32'hFFFFFFF1;
    // rom_array[45429] = 32'hFFFFFFF0;
    // rom_array[45430] = 32'hFFFFFFF0;
    // rom_array[45431] = 32'hFFFFFFF0;
    // rom_array[45432] = 32'hFFFFFFF0;
    // rom_array[45433] = 32'hFFFFFFF1;
    // rom_array[45434] = 32'hFFFFFFF1;
    // rom_array[45435] = 32'hFFFFFFF1;
    // rom_array[45436] = 32'hFFFFFFF1;
    // rom_array[45437] = 32'hFFFFFFF0;
    // rom_array[45438] = 32'hFFFFFFF0;
    // rom_array[45439] = 32'hFFFFFFF0;
    // rom_array[45440] = 32'hFFFFFFF0;
    // rom_array[45441] = 32'hFFFFFFF1;
    // rom_array[45442] = 32'hFFFFFFF1;
    // rom_array[45443] = 32'hFFFFFFF1;
    // rom_array[45444] = 32'hFFFFFFF1;
    // rom_array[45445] = 32'hFFFFFFF0;
    // rom_array[45446] = 32'hFFFFFFF0;
    // rom_array[45447] = 32'hFFFFFFF0;
    // rom_array[45448] = 32'hFFFFFFF0;
    // rom_array[45449] = 32'hFFFFFFF1;
    // rom_array[45450] = 32'hFFFFFFF1;
    // rom_array[45451] = 32'hFFFFFFF1;
    // rom_array[45452] = 32'hFFFFFFF1;
    // rom_array[45453] = 32'hFFFFFFF0;
    // rom_array[45454] = 32'hFFFFFFF0;
    // rom_array[45455] = 32'hFFFFFFF0;
    // rom_array[45456] = 32'hFFFFFFF0;
    // rom_array[45457] = 32'hFFFFFFF1;
    // rom_array[45458] = 32'hFFFFFFF1;
    // rom_array[45459] = 32'hFFFFFFF1;
    // rom_array[45460] = 32'hFFFFFFF1;
    // rom_array[45461] = 32'hFFFFFFF0;
    // rom_array[45462] = 32'hFFFFFFF0;
    // rom_array[45463] = 32'hFFFFFFF0;
    // rom_array[45464] = 32'hFFFFFFF0;
    // rom_array[45465] = 32'hFFFFFFF1;
    // rom_array[45466] = 32'hFFFFFFF1;
    // rom_array[45467] = 32'hFFFFFFF1;
    // rom_array[45468] = 32'hFFFFFFF1;
    // rom_array[45469] = 32'hFFFFFFF0;
    // rom_array[45470] = 32'hFFFFFFF0;
    // rom_array[45471] = 32'hFFFFFFF0;
    // rom_array[45472] = 32'hFFFFFFF0;
    // rom_array[45473] = 32'hFFFFFFF1;
    // rom_array[45474] = 32'hFFFFFFF1;
    // rom_array[45475] = 32'hFFFFFFF1;
    // rom_array[45476] = 32'hFFFFFFF1;
    // rom_array[45477] = 32'hFFFFFFF0;
    // rom_array[45478] = 32'hFFFFFFF0;
    // rom_array[45479] = 32'hFFFFFFF0;
    // rom_array[45480] = 32'hFFFFFFF0;
    // rom_array[45481] = 32'hFFFFFFF1;
    // rom_array[45482] = 32'hFFFFFFF1;
    // rom_array[45483] = 32'hFFFFFFF1;
    // rom_array[45484] = 32'hFFFFFFF1;
    // rom_array[45485] = 32'hFFFFFFF0;
    // rom_array[45486] = 32'hFFFFFFF0;
    // rom_array[45487] = 32'hFFFFFFF0;
    // rom_array[45488] = 32'hFFFFFFF0;
    // rom_array[45489] = 32'hFFFFFFF1;
    // rom_array[45490] = 32'hFFFFFFF1;
    // rom_array[45491] = 32'hFFFFFFF1;
    // rom_array[45492] = 32'hFFFFFFF1;
    // rom_array[45493] = 32'hFFFFFFF0;
    // rom_array[45494] = 32'hFFFFFFF0;
    // rom_array[45495] = 32'hFFFFFFF0;
    // rom_array[45496] = 32'hFFFFFFF0;
    // rom_array[45497] = 32'hFFFFFFF1;
    // rom_array[45498] = 32'hFFFFFFF1;
    // rom_array[45499] = 32'hFFFFFFF1;
    // rom_array[45500] = 32'hFFFFFFF1;
    // rom_array[45501] = 32'hFFFFFFF1;
    // rom_array[45502] = 32'hFFFFFFF1;
    // rom_array[45503] = 32'hFFFFFFF1;
    // rom_array[45504] = 32'hFFFFFFF1;
    // rom_array[45505] = 32'hFFFFFFF1;
    // rom_array[45506] = 32'hFFFFFFF1;
    // rom_array[45507] = 32'hFFFFFFF1;
    // rom_array[45508] = 32'hFFFFFFF1;
    // rom_array[45509] = 32'hFFFFFFF1;
    // rom_array[45510] = 32'hFFFFFFF1;
    // rom_array[45511] = 32'hFFFFFFF1;
    // rom_array[45512] = 32'hFFFFFFF1;
    // rom_array[45513] = 32'hFFFFFFF1;
    // rom_array[45514] = 32'hFFFFFFF1;
    // rom_array[45515] = 32'hFFFFFFF1;
    // rom_array[45516] = 32'hFFFFFFF1;
    // rom_array[45517] = 32'hFFFFFFF1;
    // rom_array[45518] = 32'hFFFFFFF1;
    // rom_array[45519] = 32'hFFFFFFF1;
    // rom_array[45520] = 32'hFFFFFFF1;
    // rom_array[45521] = 32'hFFFFFFF1;
    // rom_array[45522] = 32'hFFFFFFF1;
    // rom_array[45523] = 32'hFFFFFFF1;
    // rom_array[45524] = 32'hFFFFFFF1;
    // rom_array[45525] = 32'hFFFFFFF1;
    // rom_array[45526] = 32'hFFFFFFF1;
    // rom_array[45527] = 32'hFFFFFFF1;
    // rom_array[45528] = 32'hFFFFFFF1;
    // rom_array[45529] = 32'hFFFFFFF1;
    // rom_array[45530] = 32'hFFFFFFF1;
    // rom_array[45531] = 32'hFFFFFFF1;
    // rom_array[45532] = 32'hFFFFFFF1;
    // rom_array[45533] = 32'hFFFFFFF1;
    // rom_array[45534] = 32'hFFFFFFF1;
    // rom_array[45535] = 32'hFFFFFFF1;
    // rom_array[45536] = 32'hFFFFFFF1;
    // rom_array[45537] = 32'hFFFFFFF1;
    // rom_array[45538] = 32'hFFFFFFF1;
    // rom_array[45539] = 32'hFFFFFFF1;
    // rom_array[45540] = 32'hFFFFFFF1;
    // rom_array[45541] = 32'hFFFFFFF1;
    // rom_array[45542] = 32'hFFFFFFF1;
    // rom_array[45543] = 32'hFFFFFFF1;
    // rom_array[45544] = 32'hFFFFFFF1;
    // rom_array[45545] = 32'hFFFFFFF1;
    // rom_array[45546] = 32'hFFFFFFF1;
    // rom_array[45547] = 32'hFFFFFFF1;
    // rom_array[45548] = 32'hFFFFFFF1;
    // rom_array[45549] = 32'hFFFFFFF1;
    // rom_array[45550] = 32'hFFFFFFF1;
    // rom_array[45551] = 32'hFFFFFFF1;
    // rom_array[45552] = 32'hFFFFFFF1;
    // rom_array[45553] = 32'hFFFFFFF1;
    // rom_array[45554] = 32'hFFFFFFF1;
    // rom_array[45555] = 32'hFFFFFFF1;
    // rom_array[45556] = 32'hFFFFFFF1;
    // rom_array[45557] = 32'hFFFFFFF1;
    // rom_array[45558] = 32'hFFFFFFF1;
    // rom_array[45559] = 32'hFFFFFFF1;
    // rom_array[45560] = 32'hFFFFFFF1;
    // rom_array[45561] = 32'hFFFFFFF1;
    // rom_array[45562] = 32'hFFFFFFF1;
    // rom_array[45563] = 32'hFFFFFFF1;
    // rom_array[45564] = 32'hFFFFFFF1;
    // rom_array[45565] = 32'hFFFFFFF0;
    // rom_array[45566] = 32'hFFFFFFF0;
    // rom_array[45567] = 32'hFFFFFFF0;
    // rom_array[45568] = 32'hFFFFFFF0;
    // rom_array[45569] = 32'hFFFFFFF1;
    // rom_array[45570] = 32'hFFFFFFF1;
    // rom_array[45571] = 32'hFFFFFFF1;
    // rom_array[45572] = 32'hFFFFFFF1;
    // rom_array[45573] = 32'hFFFFFFF0;
    // rom_array[45574] = 32'hFFFFFFF0;
    // rom_array[45575] = 32'hFFFFFFF0;
    // rom_array[45576] = 32'hFFFFFFF0;
    // rom_array[45577] = 32'hFFFFFFF1;
    // rom_array[45578] = 32'hFFFFFFF1;
    // rom_array[45579] = 32'hFFFFFFF1;
    // rom_array[45580] = 32'hFFFFFFF1;
    // rom_array[45581] = 32'hFFFFFFF0;
    // rom_array[45582] = 32'hFFFFFFF0;
    // rom_array[45583] = 32'hFFFFFFF0;
    // rom_array[45584] = 32'hFFFFFFF0;
    // rom_array[45585] = 32'hFFFFFFF1;
    // rom_array[45586] = 32'hFFFFFFF1;
    // rom_array[45587] = 32'hFFFFFFF1;
    // rom_array[45588] = 32'hFFFFFFF1;
    // rom_array[45589] = 32'hFFFFFFF0;
    // rom_array[45590] = 32'hFFFFFFF0;
    // rom_array[45591] = 32'hFFFFFFF0;
    // rom_array[45592] = 32'hFFFFFFF0;
    // rom_array[45593] = 32'hFFFFFFF1;
    // rom_array[45594] = 32'hFFFFFFF1;
    // rom_array[45595] = 32'hFFFFFFF1;
    // rom_array[45596] = 32'hFFFFFFF1;
    // rom_array[45597] = 32'hFFFFFFF0;
    // rom_array[45598] = 32'hFFFFFFF0;
    // rom_array[45599] = 32'hFFFFFFF0;
    // rom_array[45600] = 32'hFFFFFFF0;
    // rom_array[45601] = 32'hFFFFFFF1;
    // rom_array[45602] = 32'hFFFFFFF1;
    // rom_array[45603] = 32'hFFFFFFF1;
    // rom_array[45604] = 32'hFFFFFFF1;
    // rom_array[45605] = 32'hFFFFFFF0;
    // rom_array[45606] = 32'hFFFFFFF0;
    // rom_array[45607] = 32'hFFFFFFF0;
    // rom_array[45608] = 32'hFFFFFFF0;
    // rom_array[45609] = 32'hFFFFFFF0;
    // rom_array[45610] = 32'hFFFFFFF0;
    // rom_array[45611] = 32'hFFFFFFF0;
    // rom_array[45612] = 32'hFFFFFFF0;
    // rom_array[45613] = 32'hFFFFFFF1;
    // rom_array[45614] = 32'hFFFFFFF1;
    // rom_array[45615] = 32'hFFFFFFF1;
    // rom_array[45616] = 32'hFFFFFFF1;
    // rom_array[45617] = 32'hFFFFFFF0;
    // rom_array[45618] = 32'hFFFFFFF0;
    // rom_array[45619] = 32'hFFFFFFF0;
    // rom_array[45620] = 32'hFFFFFFF0;
    // rom_array[45621] = 32'hFFFFFFF1;
    // rom_array[45622] = 32'hFFFFFFF1;
    // rom_array[45623] = 32'hFFFFFFF1;
    // rom_array[45624] = 32'hFFFFFFF1;
    // rom_array[45625] = 32'hFFFFFFF0;
    // rom_array[45626] = 32'hFFFFFFF0;
    // rom_array[45627] = 32'hFFFFFFF0;
    // rom_array[45628] = 32'hFFFFFFF0;
    // rom_array[45629] = 32'hFFFFFFF1;
    // rom_array[45630] = 32'hFFFFFFF1;
    // rom_array[45631] = 32'hFFFFFFF1;
    // rom_array[45632] = 32'hFFFFFFF1;
    // rom_array[45633] = 32'hFFFFFFF0;
    // rom_array[45634] = 32'hFFFFFFF0;
    // rom_array[45635] = 32'hFFFFFFF0;
    // rom_array[45636] = 32'hFFFFFFF0;
    // rom_array[45637] = 32'hFFFFFFF1;
    // rom_array[45638] = 32'hFFFFFFF1;
    // rom_array[45639] = 32'hFFFFFFF1;
    // rom_array[45640] = 32'hFFFFFFF1;
    // rom_array[45641] = 32'hFFFFFFF0;
    // rom_array[45642] = 32'hFFFFFFF0;
    // rom_array[45643] = 32'hFFFFFFF0;
    // rom_array[45644] = 32'hFFFFFFF0;
    // rom_array[45645] = 32'hFFFFFFF1;
    // rom_array[45646] = 32'hFFFFFFF1;
    // rom_array[45647] = 32'hFFFFFFF1;
    // rom_array[45648] = 32'hFFFFFFF1;
    // rom_array[45649] = 32'hFFFFFFF0;
    // rom_array[45650] = 32'hFFFFFFF0;
    // rom_array[45651] = 32'hFFFFFFF0;
    // rom_array[45652] = 32'hFFFFFFF0;
    // rom_array[45653] = 32'hFFFFFFF1;
    // rom_array[45654] = 32'hFFFFFFF1;
    // rom_array[45655] = 32'hFFFFFFF1;
    // rom_array[45656] = 32'hFFFFFFF1;
    // rom_array[45657] = 32'hFFFFFFF0;
    // rom_array[45658] = 32'hFFFFFFF0;
    // rom_array[45659] = 32'hFFFFFFF0;
    // rom_array[45660] = 32'hFFFFFFF0;
    // rom_array[45661] = 32'hFFFFFFF1;
    // rom_array[45662] = 32'hFFFFFFF1;
    // rom_array[45663] = 32'hFFFFFFF1;
    // rom_array[45664] = 32'hFFFFFFF1;
    // rom_array[45665] = 32'hFFFFFFF0;
    // rom_array[45666] = 32'hFFFFFFF0;
    // rom_array[45667] = 32'hFFFFFFF0;
    // rom_array[45668] = 32'hFFFFFFF0;
    // rom_array[45669] = 32'hFFFFFFF1;
    // rom_array[45670] = 32'hFFFFFFF1;
    // rom_array[45671] = 32'hFFFFFFF1;
    // rom_array[45672] = 32'hFFFFFFF1;
    // rom_array[45673] = 32'hFFFFFFF0;
    // rom_array[45674] = 32'hFFFFFFF0;
    // rom_array[45675] = 32'hFFFFFFF0;
    // rom_array[45676] = 32'hFFFFFFF0;
    // rom_array[45677] = 32'hFFFFFFF1;
    // rom_array[45678] = 32'hFFFFFFF1;
    // rom_array[45679] = 32'hFFFFFFF1;
    // rom_array[45680] = 32'hFFFFFFF1;
    // rom_array[45681] = 32'hFFFFFFF0;
    // rom_array[45682] = 32'hFFFFFFF0;
    // rom_array[45683] = 32'hFFFFFFF0;
    // rom_array[45684] = 32'hFFFFFFF0;
    // rom_array[45685] = 32'hFFFFFFF1;
    // rom_array[45686] = 32'hFFFFFFF1;
    // rom_array[45687] = 32'hFFFFFFF1;
    // rom_array[45688] = 32'hFFFFFFF1;
    // rom_array[45689] = 32'hFFFFFFF0;
    // rom_array[45690] = 32'hFFFFFFF0;
    // rom_array[45691] = 32'hFFFFFFF0;
    // rom_array[45692] = 32'hFFFFFFF0;
    // rom_array[45693] = 32'hFFFFFFF1;
    // rom_array[45694] = 32'hFFFFFFF1;
    // rom_array[45695] = 32'hFFFFFFF1;
    // rom_array[45696] = 32'hFFFFFFF1;
    // rom_array[45697] = 32'hFFFFFFF0;
    // rom_array[45698] = 32'hFFFFFFF0;
    // rom_array[45699] = 32'hFFFFFFF0;
    // rom_array[45700] = 32'hFFFFFFF0;
    // rom_array[45701] = 32'hFFFFFFF1;
    // rom_array[45702] = 32'hFFFFFFF1;
    // rom_array[45703] = 32'hFFFFFFF1;
    // rom_array[45704] = 32'hFFFFFFF1;
    // rom_array[45705] = 32'hFFFFFFF0;
    // rom_array[45706] = 32'hFFFFFFF0;
    // rom_array[45707] = 32'hFFFFFFF0;
    // rom_array[45708] = 32'hFFFFFFF0;
    // rom_array[45709] = 32'hFFFFFFF1;
    // rom_array[45710] = 32'hFFFFFFF1;
    // rom_array[45711] = 32'hFFFFFFF1;
    // rom_array[45712] = 32'hFFFFFFF1;
    // rom_array[45713] = 32'hFFFFFFF0;
    // rom_array[45714] = 32'hFFFFFFF0;
    // rom_array[45715] = 32'hFFFFFFF0;
    // rom_array[45716] = 32'hFFFFFFF0;
    // rom_array[45717] = 32'hFFFFFFF1;
    // rom_array[45718] = 32'hFFFFFFF1;
    // rom_array[45719] = 32'hFFFFFFF1;
    // rom_array[45720] = 32'hFFFFFFF1;
    // rom_array[45721] = 32'hFFFFFFF0;
    // rom_array[45722] = 32'hFFFFFFF0;
    // rom_array[45723] = 32'hFFFFFFF0;
    // rom_array[45724] = 32'hFFFFFFF0;
    // rom_array[45725] = 32'hFFFFFFF1;
    // rom_array[45726] = 32'hFFFFFFF1;
    // rom_array[45727] = 32'hFFFFFFF1;
    // rom_array[45728] = 32'hFFFFFFF1;
    // rom_array[45729] = 32'hFFFFFFF0;
    // rom_array[45730] = 32'hFFFFFFF0;
    // rom_array[45731] = 32'hFFFFFFF0;
    // rom_array[45732] = 32'hFFFFFFF0;
    // rom_array[45733] = 32'hFFFFFFF1;
    // rom_array[45734] = 32'hFFFFFFF1;
    // rom_array[45735] = 32'hFFFFFFF1;
    // rom_array[45736] = 32'hFFFFFFF1;
    // rom_array[45737] = 32'hFFFFFFF0;
    // rom_array[45738] = 32'hFFFFFFF0;
    // rom_array[45739] = 32'hFFFFFFF0;
    // rom_array[45740] = 32'hFFFFFFF0;
    // rom_array[45741] = 32'hFFFFFFF1;
    // rom_array[45742] = 32'hFFFFFFF1;
    // rom_array[45743] = 32'hFFFFFFF1;
    // rom_array[45744] = 32'hFFFFFFF1;
    // rom_array[45745] = 32'hFFFFFFF0;
    // rom_array[45746] = 32'hFFFFFFF0;
    // rom_array[45747] = 32'hFFFFFFF0;
    // rom_array[45748] = 32'hFFFFFFF0;
    // rom_array[45749] = 32'hFFFFFFF1;
    // rom_array[45750] = 32'hFFFFFFF1;
    // rom_array[45751] = 32'hFFFFFFF1;
    // rom_array[45752] = 32'hFFFFFFF1;
    // rom_array[45753] = 32'hFFFFFFF0;
    // rom_array[45754] = 32'hFFFFFFF0;
    // rom_array[45755] = 32'hFFFFFFF0;
    // rom_array[45756] = 32'hFFFFFFF0;
    // rom_array[45757] = 32'hFFFFFFF1;
    // rom_array[45758] = 32'hFFFFFFF1;
    // rom_array[45759] = 32'hFFFFFFF1;
    // rom_array[45760] = 32'hFFFFFFF1;
    // rom_array[45761] = 32'hFFFFFFF0;
    // rom_array[45762] = 32'hFFFFFFF0;
    // rom_array[45763] = 32'hFFFFFFF0;
    // rom_array[45764] = 32'hFFFFFFF0;
    // rom_array[45765] = 32'hFFFFFFF1;
    // rom_array[45766] = 32'hFFFFFFF1;
    // rom_array[45767] = 32'hFFFFFFF1;
    // rom_array[45768] = 32'hFFFFFFF1;
    // rom_array[45769] = 32'hFFFFFFF0;
    // rom_array[45770] = 32'hFFFFFFF0;
    // rom_array[45771] = 32'hFFFFFFF0;
    // rom_array[45772] = 32'hFFFFFFF0;
    // rom_array[45773] = 32'hFFFFFFF1;
    // rom_array[45774] = 32'hFFFFFFF1;
    // rom_array[45775] = 32'hFFFFFFF1;
    // rom_array[45776] = 32'hFFFFFFF1;
    // rom_array[45777] = 32'hFFFFFFF0;
    // rom_array[45778] = 32'hFFFFFFF0;
    // rom_array[45779] = 32'hFFFFFFF0;
    // rom_array[45780] = 32'hFFFFFFF0;
    // rom_array[45781] = 32'hFFFFFFF1;
    // rom_array[45782] = 32'hFFFFFFF1;
    // rom_array[45783] = 32'hFFFFFFF1;
    // rom_array[45784] = 32'hFFFFFFF1;
    // rom_array[45785] = 32'hFFFFFFF1;
    // rom_array[45786] = 32'hFFFFFFF1;
    // rom_array[45787] = 32'hFFFFFFF1;
    // rom_array[45788] = 32'hFFFFFFF1;
    // rom_array[45789] = 32'hFFFFFFF1;
    // rom_array[45790] = 32'hFFFFFFF1;
    // rom_array[45791] = 32'hFFFFFFF1;
    // rom_array[45792] = 32'hFFFFFFF1;
    // rom_array[45793] = 32'hFFFFFFF1;
    // rom_array[45794] = 32'hFFFFFFF1;
    // rom_array[45795] = 32'hFFFFFFF1;
    // rom_array[45796] = 32'hFFFFFFF1;
    // rom_array[45797] = 32'hFFFFFFF1;
    // rom_array[45798] = 32'hFFFFFFF1;
    // rom_array[45799] = 32'hFFFFFFF1;
    // rom_array[45800] = 32'hFFFFFFF1;
    // rom_array[45801] = 32'hFFFFFFF1;
    // rom_array[45802] = 32'hFFFFFFF1;
    // rom_array[45803] = 32'hFFFFFFF1;
    // rom_array[45804] = 32'hFFFFFFF1;
    // rom_array[45805] = 32'hFFFFFFF1;
    // rom_array[45806] = 32'hFFFFFFF1;
    // rom_array[45807] = 32'hFFFFFFF1;
    // rom_array[45808] = 32'hFFFFFFF1;
    // rom_array[45809] = 32'hFFFFFFF1;
    // rom_array[45810] = 32'hFFFFFFF1;
    // rom_array[45811] = 32'hFFFFFFF1;
    // rom_array[45812] = 32'hFFFFFFF1;
    // rom_array[45813] = 32'hFFFFFFF1;
    // rom_array[45814] = 32'hFFFFFFF1;
    // rom_array[45815] = 32'hFFFFFFF1;
    // rom_array[45816] = 32'hFFFFFFF1;
    // rom_array[45817] = 32'hFFFFFFF1;
    // rom_array[45818] = 32'hFFFFFFF1;
    // rom_array[45819] = 32'hFFFFFFF1;
    // rom_array[45820] = 32'hFFFFFFF1;
    // rom_array[45821] = 32'hFFFFFFF1;
    // rom_array[45822] = 32'hFFFFFFF1;
    // rom_array[45823] = 32'hFFFFFFF1;
    // rom_array[45824] = 32'hFFFFFFF1;
    // rom_array[45825] = 32'hFFFFFFF1;
    // rom_array[45826] = 32'hFFFFFFF1;
    // rom_array[45827] = 32'hFFFFFFF1;
    // rom_array[45828] = 32'hFFFFFFF1;
    // rom_array[45829] = 32'hFFFFFFF1;
    // rom_array[45830] = 32'hFFFFFFF1;
    // rom_array[45831] = 32'hFFFFFFF1;
    // rom_array[45832] = 32'hFFFFFFF1;
    // rom_array[45833] = 32'hFFFFFFF1;
    // rom_array[45834] = 32'hFFFFFFF1;
    // rom_array[45835] = 32'hFFFFFFF1;
    // rom_array[45836] = 32'hFFFFFFF1;
    // rom_array[45837] = 32'hFFFFFFF0;
    // rom_array[45838] = 32'hFFFFFFF0;
    // rom_array[45839] = 32'hFFFFFFF0;
    // rom_array[45840] = 32'hFFFFFFF0;
    // rom_array[45841] = 32'hFFFFFFF1;
    // rom_array[45842] = 32'hFFFFFFF1;
    // rom_array[45843] = 32'hFFFFFFF1;
    // rom_array[45844] = 32'hFFFFFFF1;
    // rom_array[45845] = 32'hFFFFFFF0;
    // rom_array[45846] = 32'hFFFFFFF0;
    // rom_array[45847] = 32'hFFFFFFF0;
    // rom_array[45848] = 32'hFFFFFFF0;
    // rom_array[45849] = 32'hFFFFFFF1;
    // rom_array[45850] = 32'hFFFFFFF1;
    // rom_array[45851] = 32'hFFFFFFF1;
    // rom_array[45852] = 32'hFFFFFFF1;
    // rom_array[45853] = 32'hFFFFFFF0;
    // rom_array[45854] = 32'hFFFFFFF0;
    // rom_array[45855] = 32'hFFFFFFF0;
    // rom_array[45856] = 32'hFFFFFFF0;
    // rom_array[45857] = 32'hFFFFFFF1;
    // rom_array[45858] = 32'hFFFFFFF1;
    // rom_array[45859] = 32'hFFFFFFF1;
    // rom_array[45860] = 32'hFFFFFFF1;
    // rom_array[45861] = 32'hFFFFFFF0;
    // rom_array[45862] = 32'hFFFFFFF0;
    // rom_array[45863] = 32'hFFFFFFF0;
    // rom_array[45864] = 32'hFFFFFFF0;
    // rom_array[45865] = 32'hFFFFFFF1;
    // rom_array[45866] = 32'hFFFFFFF1;
    // rom_array[45867] = 32'hFFFFFFF1;
    // rom_array[45868] = 32'hFFFFFFF1;
    // rom_array[45869] = 32'hFFFFFFF0;
    // rom_array[45870] = 32'hFFFFFFF0;
    // rom_array[45871] = 32'hFFFFFFF0;
    // rom_array[45872] = 32'hFFFFFFF0;
    // rom_array[45873] = 32'hFFFFFFF1;
    // rom_array[45874] = 32'hFFFFFFF1;
    // rom_array[45875] = 32'hFFFFFFF1;
    // rom_array[45876] = 32'hFFFFFFF1;
    // rom_array[45877] = 32'hFFFFFFF0;
    // rom_array[45878] = 32'hFFFFFFF0;
    // rom_array[45879] = 32'hFFFFFFF0;
    // rom_array[45880] = 32'hFFFFFFF0;
    // rom_array[45881] = 32'hFFFFFFF1;
    // rom_array[45882] = 32'hFFFFFFF1;
    // rom_array[45883] = 32'hFFFFFFF1;
    // rom_array[45884] = 32'hFFFFFFF1;
    // rom_array[45885] = 32'hFFFFFFF0;
    // rom_array[45886] = 32'hFFFFFFF0;
    // rom_array[45887] = 32'hFFFFFFF0;
    // rom_array[45888] = 32'hFFFFFFF0;
    // rom_array[45889] = 32'hFFFFFFF1;
    // rom_array[45890] = 32'hFFFFFFF1;
    // rom_array[45891] = 32'hFFFFFFF1;
    // rom_array[45892] = 32'hFFFFFFF1;
    // rom_array[45893] = 32'hFFFFFFF0;
    // rom_array[45894] = 32'hFFFFFFF0;
    // rom_array[45895] = 32'hFFFFFFF0;
    // rom_array[45896] = 32'hFFFFFFF0;
    // rom_array[45897] = 32'hFFFFFFF1;
    // rom_array[45898] = 32'hFFFFFFF1;
    // rom_array[45899] = 32'hFFFFFFF1;
    // rom_array[45900] = 32'hFFFFFFF1;
    // rom_array[45901] = 32'hFFFFFFF0;
    // rom_array[45902] = 32'hFFFFFFF0;
    // rom_array[45903] = 32'hFFFFFFF0;
    // rom_array[45904] = 32'hFFFFFFF0;
    // rom_array[45905] = 32'hFFFFFFF1;
    // rom_array[45906] = 32'hFFFFFFF1;
    // rom_array[45907] = 32'hFFFFFFF1;
    // rom_array[45908] = 32'hFFFFFFF1;
    // rom_array[45909] = 32'hFFFFFFF0;
    // rom_array[45910] = 32'hFFFFFFF0;
    // rom_array[45911] = 32'hFFFFFFF0;
    // rom_array[45912] = 32'hFFFFFFF0;
    // rom_array[45913] = 32'hFFFFFFF1;
    // rom_array[45914] = 32'hFFFFFFF1;
    // rom_array[45915] = 32'hFFFFFFF1;
    // rom_array[45916] = 32'hFFFFFFF1;
    // rom_array[45917] = 32'hFFFFFFF0;
    // rom_array[45918] = 32'hFFFFFFF0;
    // rom_array[45919] = 32'hFFFFFFF0;
    // rom_array[45920] = 32'hFFFFFFF0;
    // rom_array[45921] = 32'hFFFFFFF1;
    // rom_array[45922] = 32'hFFFFFFF1;
    // rom_array[45923] = 32'hFFFFFFF1;
    // rom_array[45924] = 32'hFFFFFFF1;
    // rom_array[45925] = 32'hFFFFFFF0;
    // rom_array[45926] = 32'hFFFFFFF0;
    // rom_array[45927] = 32'hFFFFFFF0;
    // rom_array[45928] = 32'hFFFFFFF0;
    // rom_array[45929] = 32'hFFFFFFF1;
    // rom_array[45930] = 32'hFFFFFFF1;
    // rom_array[45931] = 32'hFFFFFFF1;
    // rom_array[45932] = 32'hFFFFFFF1;
    // rom_array[45933] = 32'hFFFFFFF0;
    // rom_array[45934] = 32'hFFFFFFF0;
    // rom_array[45935] = 32'hFFFFFFF0;
    // rom_array[45936] = 32'hFFFFFFF0;
    // rom_array[45937] = 32'hFFFFFFF1;
    // rom_array[45938] = 32'hFFFFFFF1;
    // rom_array[45939] = 32'hFFFFFFF1;
    // rom_array[45940] = 32'hFFFFFFF1;
    // rom_array[45941] = 32'hFFFFFFF0;
    // rom_array[45942] = 32'hFFFFFFF0;
    // rom_array[45943] = 32'hFFFFFFF0;
    // rom_array[45944] = 32'hFFFFFFF0;
    // rom_array[45945] = 32'hFFFFFFF1;
    // rom_array[45946] = 32'hFFFFFFF1;
    // rom_array[45947] = 32'hFFFFFFF1;
    // rom_array[45948] = 32'hFFFFFFF1;
    // rom_array[45949] = 32'hFFFFFFF0;
    // rom_array[45950] = 32'hFFFFFFF0;
    // rom_array[45951] = 32'hFFFFFFF0;
    // rom_array[45952] = 32'hFFFFFFF0;
    // rom_array[45953] = 32'hFFFFFFF1;
    // rom_array[45954] = 32'hFFFFFFF1;
    // rom_array[45955] = 32'hFFFFFFF1;
    // rom_array[45956] = 32'hFFFFFFF1;
    // rom_array[45957] = 32'hFFFFFFF0;
    // rom_array[45958] = 32'hFFFFFFF0;
    // rom_array[45959] = 32'hFFFFFFF0;
    // rom_array[45960] = 32'hFFFFFFF0;
    // rom_array[45961] = 32'hFFFFFFF1;
    // rom_array[45962] = 32'hFFFFFFF1;
    // rom_array[45963] = 32'hFFFFFFF1;
    // rom_array[45964] = 32'hFFFFFFF1;
    // rom_array[45965] = 32'hFFFFFFF0;
    // rom_array[45966] = 32'hFFFFFFF0;
    // rom_array[45967] = 32'hFFFFFFF0;
    // rom_array[45968] = 32'hFFFFFFF0;
    // rom_array[45969] = 32'hFFFFFFF1;
    // rom_array[45970] = 32'hFFFFFFF1;
    // rom_array[45971] = 32'hFFFFFFF1;
    // rom_array[45972] = 32'hFFFFFFF1;
    // rom_array[45973] = 32'hFFFFFFF0;
    // rom_array[45974] = 32'hFFFFFFF0;
    // rom_array[45975] = 32'hFFFFFFF0;
    // rom_array[45976] = 32'hFFFFFFF0;
    // rom_array[45977] = 32'hFFFFFFF1;
    // rom_array[45978] = 32'hFFFFFFF1;
    // rom_array[45979] = 32'hFFFFFFF1;
    // rom_array[45980] = 32'hFFFFFFF1;
    // rom_array[45981] = 32'hFFFFFFF0;
    // rom_array[45982] = 32'hFFFFFFF0;
    // rom_array[45983] = 32'hFFFFFFF0;
    // rom_array[45984] = 32'hFFFFFFF0;
    // rom_array[45985] = 32'hFFFFFFF1;
    // rom_array[45986] = 32'hFFFFFFF1;
    // rom_array[45987] = 32'hFFFFFFF1;
    // rom_array[45988] = 32'hFFFFFFF1;
    // rom_array[45989] = 32'hFFFFFFF0;
    // rom_array[45990] = 32'hFFFFFFF0;
    // rom_array[45991] = 32'hFFFFFFF0;
    // rom_array[45992] = 32'hFFFFFFF0;
    // rom_array[45993] = 32'hFFFFFFF1;
    // rom_array[45994] = 32'hFFFFFFF1;
    // rom_array[45995] = 32'hFFFFFFF1;
    // rom_array[45996] = 32'hFFFFFFF1;
    // rom_array[45997] = 32'hFFFFFFF0;
    // rom_array[45998] = 32'hFFFFFFF0;
    // rom_array[45999] = 32'hFFFFFFF0;
    // rom_array[46000] = 32'hFFFFFFF0;
    // rom_array[46001] = 32'hFFFFFFF1;
    // rom_array[46002] = 32'hFFFFFFF1;
    // rom_array[46003] = 32'hFFFFFFF1;
    // rom_array[46004] = 32'hFFFFFFF1;
    // rom_array[46005] = 32'hFFFFFFF0;
    // rom_array[46006] = 32'hFFFFFFF0;
    // rom_array[46007] = 32'hFFFFFFF0;
    // rom_array[46008] = 32'hFFFFFFF0;


end

always_ff @(posedge clk) begin
    if(ren1 || ren2) begin
        dout1 <= rom_array[addr1];
        dout2 <= rom_array[addr2];
    end
end

endmodule
